//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: bram]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- BEGIN Grid Verilog module: grid_bram -----
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for grid_bram -----
module grid_bram(global_resetn,
                 scan_en,
                 scan_mode,
                 top_width_0_height_0_subtile_0__pin_I00_0_,
                 top_width_0_height_0_subtile_0__pin_I00_1_,
                 top_width_0_height_0_subtile_0__pin_I00_2_,
                 top_width_0_height_0_subtile_0__pin_I00_3_,
                 top_width_0_height_0_subtile_0__pin_I00_4_,
                 top_width_0_height_0_subtile_0__pin_I00_5_,
                 top_width_0_height_0_subtile_0__pin_I00_6_,
                 top_width_0_height_0_subtile_0__pin_I00_7_,
                 top_width_0_height_0_subtile_0__pin_I00_8_,
                 top_width_0_height_0_subtile_0__pin_I00_9_,
                 top_width_0_height_0_subtile_0__pin_I00_10_,
                 top_width_0_height_0_subtile_0__pin_I00_11_,
                 top_width_0_height_0_subtile_0__pin_I10_0_,
                 top_width_0_height_0_subtile_0__pin_I10_1_,
                 top_width_0_height_0_subtile_0__pin_I10_2_,
                 top_width_0_height_0_subtile_0__pin_I10_3_,
                 top_width_0_height_0_subtile_0__pin_I10_4_,
                 top_width_0_height_0_subtile_0__pin_I10_5_,
                 top_width_0_height_0_subtile_0__pin_I10_6_,
                 top_width_0_height_0_subtile_0__pin_I10_7_,
                 top_width_0_height_0_subtile_0__pin_I10_8_,
                 top_width_0_height_0_subtile_0__pin_I10_9_,
                 top_width_0_height_0_subtile_0__pin_I10_10_,
                 top_width_0_height_0_subtile_0__pin_I10_11_,
                 top_width_0_height_0_subtile_0__pin_IS0_0_,
                 top_width_0_height_0_subtile_0__pin_IS0_1_,
                 top_width_0_height_0_subtile_0__pin_IS0_2_,
                 top_width_0_height_1_subtile_0__pin_I01_0_,
                 top_width_0_height_1_subtile_0__pin_I01_1_,
                 top_width_0_height_1_subtile_0__pin_I01_2_,
                 top_width_0_height_1_subtile_0__pin_I01_3_,
                 top_width_0_height_1_subtile_0__pin_I01_4_,
                 top_width_0_height_1_subtile_0__pin_I01_5_,
                 top_width_0_height_1_subtile_0__pin_I01_6_,
                 top_width_0_height_1_subtile_0__pin_I01_7_,
                 top_width_0_height_1_subtile_0__pin_I01_8_,
                 top_width_0_height_1_subtile_0__pin_I01_9_,
                 top_width_0_height_1_subtile_0__pin_I01_10_,
                 top_width_0_height_1_subtile_0__pin_I01_11_,
                 top_width_0_height_1_subtile_0__pin_I11_0_,
                 top_width_0_height_1_subtile_0__pin_I11_1_,
                 top_width_0_height_1_subtile_0__pin_I11_2_,
                 top_width_0_height_1_subtile_0__pin_I11_3_,
                 top_width_0_height_1_subtile_0__pin_I11_4_,
                 top_width_0_height_1_subtile_0__pin_I11_5_,
                 top_width_0_height_1_subtile_0__pin_I11_6_,
                 top_width_0_height_1_subtile_0__pin_I11_7_,
                 top_width_0_height_1_subtile_0__pin_I11_8_,
                 top_width_0_height_1_subtile_0__pin_I11_9_,
                 top_width_0_height_1_subtile_0__pin_I11_10_,
                 top_width_0_height_1_subtile_0__pin_I11_11_,
                 top_width_0_height_1_subtile_0__pin_IS1_0_,
                 top_width_0_height_1_subtile_0__pin_IS1_1_,
                 top_width_0_height_1_subtile_0__pin_IS1_2_,
                 top_width_0_height_2_subtile_0__pin_I02_0_,
                 top_width_0_height_2_subtile_0__pin_I02_1_,
                 top_width_0_height_2_subtile_0__pin_I02_2_,
                 top_width_0_height_2_subtile_0__pin_I02_3_,
                 top_width_0_height_2_subtile_0__pin_I02_4_,
                 top_width_0_height_2_subtile_0__pin_I02_5_,
                 top_width_0_height_2_subtile_0__pin_I02_6_,
                 top_width_0_height_2_subtile_0__pin_I02_7_,
                 top_width_0_height_2_subtile_0__pin_I02_8_,
                 top_width_0_height_2_subtile_0__pin_I02_9_,
                 top_width_0_height_2_subtile_0__pin_I02_10_,
                 top_width_0_height_2_subtile_0__pin_I02_11_,
                 top_width_0_height_2_subtile_0__pin_I12_0_,
                 top_width_0_height_2_subtile_0__pin_I12_1_,
                 top_width_0_height_2_subtile_0__pin_I12_2_,
                 top_width_0_height_2_subtile_0__pin_I12_3_,
                 top_width_0_height_2_subtile_0__pin_I12_4_,
                 top_width_0_height_2_subtile_0__pin_I12_5_,
                 top_width_0_height_2_subtile_0__pin_I12_6_,
                 top_width_0_height_2_subtile_0__pin_I12_7_,
                 top_width_0_height_2_subtile_0__pin_I12_8_,
                 top_width_0_height_2_subtile_0__pin_I12_9_,
                 top_width_0_height_2_subtile_0__pin_I12_10_,
                 top_width_0_height_2_subtile_0__pin_I12_11_,
                 top_width_0_height_2_subtile_0__pin_IS2_0_,
                 top_width_0_height_2_subtile_0__pin_IS2_1_,
                 top_width_0_height_2_subtile_0__pin_IS2_2_,
                 top_width_0_height_2_subtile_0__pin_PL_INIT_i_0_,
                 top_width_0_height_2_subtile_0__pin_PL_ENA_i_0_,
                 top_width_0_height_2_subtile_0__pin_PL_REN_i_0_,
                 top_width_0_height_2_subtile_0__pin_PL_WEN_i_0_,
                 top_width_0_height_2_subtile_0__pin_PL_WEN_i_1_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_0_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_1_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_2_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_3_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_4_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_5_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_6_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_7_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_8_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_9_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_10_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_11_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_12_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_13_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_14_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_15_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_16_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_17_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_18_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_19_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_20_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_21_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_22_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_23_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_24_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_25_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_26_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_27_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_28_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_29_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_30_,
                 top_width_0_height_2_subtile_0__pin_PL_ADDR_i_31_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_0_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_1_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_2_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_3_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_4_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_5_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_6_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_7_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_8_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_9_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_10_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_11_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_12_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_13_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_14_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_15_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_16_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_17_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_18_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_19_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_20_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_21_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_22_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_23_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_24_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_25_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_26_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_27_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_28_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_29_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_30_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_31_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_32_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_33_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_34_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_i_35_,
                 top_width_0_height_2_subtile_0__pin_PL_CLK_i_0_,
                 right_width_0_height_0_subtile_0__pin_I20_0_,
                 right_width_0_height_0_subtile_0__pin_I20_1_,
                 right_width_0_height_0_subtile_0__pin_I20_2_,
                 right_width_0_height_0_subtile_0__pin_I20_3_,
                 right_width_0_height_0_subtile_0__pin_I20_4_,
                 right_width_0_height_0_subtile_0__pin_I20_5_,
                 right_width_0_height_0_subtile_0__pin_I20_6_,
                 right_width_0_height_0_subtile_0__pin_I20_7_,
                 right_width_0_height_0_subtile_0__pin_I20_8_,
                 right_width_0_height_0_subtile_0__pin_I20_9_,
                 right_width_0_height_0_subtile_0__pin_I20_10_,
                 right_width_0_height_0_subtile_0__pin_I20_11_,
                 right_width_0_height_0_subtile_0__pin_I30_0_,
                 right_width_0_height_0_subtile_0__pin_I30_1_,
                 right_width_0_height_0_subtile_0__pin_I30_2_,
                 right_width_0_height_0_subtile_0__pin_I30_3_,
                 right_width_0_height_0_subtile_0__pin_I30_4_,
                 right_width_0_height_0_subtile_0__pin_I30_5_,
                 right_width_0_height_0_subtile_0__pin_I30_6_,
                 right_width_0_height_0_subtile_0__pin_I30_7_,
                 right_width_0_height_0_subtile_0__pin_I30_8_,
                 right_width_0_height_0_subtile_0__pin_I30_9_,
                 right_width_0_height_0_subtile_0__pin_I30_10_,
                 right_width_0_height_0_subtile_0__pin_I30_11_,
                 right_width_0_height_0_subtile_0__pin_IS0_3_,
                 right_width_0_height_0_subtile_0__pin_IS0_4_,
                 right_width_0_height_0_subtile_0__pin_IS0_5_,
                 right_width_0_height_0_subtile_0__pin_sr_in_0_,
                 right_width_0_height_0_subtile_0__pin_sr_in_1_,
                 right_width_0_height_0_subtile_0__pin_sr_in_2_,
                 right_width_0_height_0_subtile_0__pin_sr_in_3_,
                 right_width_0_height_0_subtile_0__pin_sr_in_4_,
                 right_width_0_height_0_subtile_0__pin_sr_in_5_,
                 right_width_0_height_0_subtile_0__pin_plr_i_0_,
                 right_width_0_height_0_subtile_0__pin_plr_i_1_,
                 right_width_0_height_0_subtile_0__pin_plr_i_2_,
                 right_width_0_height_0_subtile_0__pin_plr_i_3_,
                 right_width_0_height_0_subtile_0__pin_plr_i_4_,
                 right_width_0_height_0_subtile_0__pin_plr_i_5_,
                 right_width_0_height_0_subtile_0__pin_plr_i_6_,
                 right_width_0_height_0_subtile_0__pin_plr_i_7_,
                 right_width_0_height_0_subtile_0__pin_plr_i_8_,
                 right_width_0_height_0_subtile_0__pin_plr_i_9_,
                 right_width_0_height_0_subtile_0__pin_plr_i_10_,
                 right_width_0_height_0_subtile_0__pin_plr_i_11_,
                 right_width_0_height_0_subtile_0__pin_plr_i_12_,
                 right_width_0_height_0_subtile_0__pin_plr_i_13_,
                 right_width_0_height_0_subtile_0__pin_plr_i_14_,
                 right_width_0_height_0_subtile_0__pin_plr_i_15_,
                 right_width_0_height_0_subtile_0__pin_plr_i_16_,
                 right_width_0_height_0_subtile_0__pin_plr_i_17_,
                 right_width_0_height_0_subtile_0__pin_plr_i_18_,
                 right_width_0_height_0_subtile_0__pin_plr_i_19_,
                 right_width_0_height_0_subtile_0__pin_plr_i_20_,
                 right_width_0_height_0_subtile_0__pin_plr_i_21_,
                 right_width_0_height_0_subtile_0__pin_plr_i_22_,
                 right_width_0_height_0_subtile_0__pin_plr_i_23_,
                 right_width_0_height_0_subtile_0__pin_plr_i_24_,
                 right_width_0_height_0_subtile_0__pin_plr_i_25_,
                 right_width_0_height_0_subtile_0__pin_plr_i_26_,
                 right_width_0_height_0_subtile_0__pin_plr_i_27_,
                 right_width_0_height_0_subtile_0__pin_plr_i_28_,
                 right_width_0_height_0_subtile_0__pin_plr_i_29_,
                 right_width_0_height_0_subtile_0__pin_plr_i_30_,
                 right_width_0_height_0_subtile_0__pin_plr_i_31_,
                 right_width_0_height_0_subtile_0__pin_plr_i_32_,
                 right_width_0_height_0_subtile_0__pin_plr_i_33_,
                 right_width_0_height_0_subtile_0__pin_plr_i_34_,
                 right_width_0_height_0_subtile_0__pin_plr_i_35_,
                 right_width_0_height_1_subtile_0__pin_I21_0_,
                 right_width_0_height_1_subtile_0__pin_I21_1_,
                 right_width_0_height_1_subtile_0__pin_I21_2_,
                 right_width_0_height_1_subtile_0__pin_I21_3_,
                 right_width_0_height_1_subtile_0__pin_I21_4_,
                 right_width_0_height_1_subtile_0__pin_I21_5_,
                 right_width_0_height_1_subtile_0__pin_I21_6_,
                 right_width_0_height_1_subtile_0__pin_I21_7_,
                 right_width_0_height_1_subtile_0__pin_I21_8_,
                 right_width_0_height_1_subtile_0__pin_I21_9_,
                 right_width_0_height_1_subtile_0__pin_I21_10_,
                 right_width_0_height_1_subtile_0__pin_I21_11_,
                 right_width_0_height_1_subtile_0__pin_I31_0_,
                 right_width_0_height_1_subtile_0__pin_I31_1_,
                 right_width_0_height_1_subtile_0__pin_I31_2_,
                 right_width_0_height_1_subtile_0__pin_I31_3_,
                 right_width_0_height_1_subtile_0__pin_I31_4_,
                 right_width_0_height_1_subtile_0__pin_I31_5_,
                 right_width_0_height_1_subtile_0__pin_I31_6_,
                 right_width_0_height_1_subtile_0__pin_I31_7_,
                 right_width_0_height_1_subtile_0__pin_I31_8_,
                 right_width_0_height_1_subtile_0__pin_I31_9_,
                 right_width_0_height_1_subtile_0__pin_I31_10_,
                 right_width_0_height_1_subtile_0__pin_I31_11_,
                 right_width_0_height_1_subtile_0__pin_IS1_3_,
                 right_width_0_height_1_subtile_0__pin_IS1_4_,
                 right_width_0_height_1_subtile_0__pin_IS1_5_,
                 right_width_0_height_2_subtile_0__pin_I22_0_,
                 right_width_0_height_2_subtile_0__pin_I22_1_,
                 right_width_0_height_2_subtile_0__pin_I22_2_,
                 right_width_0_height_2_subtile_0__pin_I22_3_,
                 right_width_0_height_2_subtile_0__pin_I22_4_,
                 right_width_0_height_2_subtile_0__pin_I22_5_,
                 right_width_0_height_2_subtile_0__pin_I22_6_,
                 right_width_0_height_2_subtile_0__pin_I22_7_,
                 right_width_0_height_2_subtile_0__pin_I22_8_,
                 right_width_0_height_2_subtile_0__pin_I22_9_,
                 right_width_0_height_2_subtile_0__pin_I22_10_,
                 right_width_0_height_2_subtile_0__pin_I22_11_,
                 right_width_0_height_2_subtile_0__pin_I32_0_,
                 right_width_0_height_2_subtile_0__pin_I32_1_,
                 right_width_0_height_2_subtile_0__pin_I32_2_,
                 right_width_0_height_2_subtile_0__pin_I32_3_,
                 right_width_0_height_2_subtile_0__pin_I32_4_,
                 right_width_0_height_2_subtile_0__pin_I32_5_,
                 right_width_0_height_2_subtile_0__pin_I32_6_,
                 right_width_0_height_2_subtile_0__pin_I32_7_,
                 right_width_0_height_2_subtile_0__pin_I32_8_,
                 right_width_0_height_2_subtile_0__pin_I32_9_,
                 right_width_0_height_2_subtile_0__pin_I32_10_,
                 right_width_0_height_2_subtile_0__pin_I32_11_,
                 right_width_0_height_2_subtile_0__pin_IS2_3_,
                 right_width_0_height_2_subtile_0__pin_IS2_4_,
                 right_width_0_height_2_subtile_0__pin_IS2_5_,
                 left_width_0_height_0_subtile_0__pin_sc_in_0_,
                 left_width_0_height_0_subtile_0__pin_sc_in_1_,
                 left_width_0_height_0_subtile_0__pin_sc_in_2_,
                 left_width_0_height_0_subtile_0__pin_sc_in_3_,
                 left_width_0_height_0_subtile_0__pin_sc_in_4_,
                 left_width_0_height_0_subtile_0__pin_sc_in_5_,
                 left_width_0_height_0_subtile_0__pin_clk_0_,
                 left_width_0_height_0_subtile_0__pin_clk_1_,
                 left_width_0_height_0_subtile_0__pin_clk_2_,
                 left_width_0_height_0_subtile_0__pin_clk_3_,
                 left_width_0_height_0_subtile_0__pin_clk_4_,
                 left_width_0_height_0_subtile_0__pin_clk_5_,
                 left_width_0_height_0_subtile_0__pin_clk_6_,
                 left_width_0_height_0_subtile_0__pin_clk_7_,
                 left_width_0_height_0_subtile_0__pin_clk_8_,
                 left_width_0_height_0_subtile_0__pin_clk_9_,
                 left_width_0_height_0_subtile_0__pin_clk_10_,
                 left_width_0_height_0_subtile_0__pin_clk_11_,
                 left_width_0_height_0_subtile_0__pin_clk_12_,
                 left_width_0_height_0_subtile_0__pin_clk_13_,
                 left_width_0_height_0_subtile_0__pin_clk_14_,
                 left_width_0_height_0_subtile_0__pin_clk_15_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_0_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_1_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_2_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_3_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_4_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_5_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_6_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_7_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_8_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_9_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_10_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_11_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_12_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_13_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_14_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_15_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_16_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_17_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_18_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_19_,
                 bl,
                 wl,
                 top_width_0_height_0_subtile_0__pin_O0_0_,
                 top_width_0_height_0_subtile_0__pin_O0_1_,
                 top_width_0_height_0_subtile_0__pin_O0_2_,
                 top_width_0_height_0_subtile_0__pin_O0_3_,
                 top_width_0_height_0_subtile_0__pin_O0_4_,
                 top_width_0_height_0_subtile_0__pin_O0_5_,
                 top_width_0_height_0_subtile_0__pin_O0_6_,
                 top_width_0_height_0_subtile_0__pin_O0_7_,
                 top_width_0_height_0_subtile_0__pin_O0_8_,
                 top_width_0_height_0_subtile_0__pin_O0_9_,
                 top_width_0_height_0_subtile_0__pin_O0_10_,
                 top_width_0_height_0_subtile_0__pin_O0_11_,
                 top_width_0_height_1_subtile_0__pin_O1_0_,
                 top_width_0_height_1_subtile_0__pin_O1_1_,
                 top_width_0_height_1_subtile_0__pin_O1_2_,
                 top_width_0_height_1_subtile_0__pin_O1_3_,
                 top_width_0_height_1_subtile_0__pin_O1_4_,
                 top_width_0_height_1_subtile_0__pin_O1_5_,
                 top_width_0_height_1_subtile_0__pin_O1_6_,
                 top_width_0_height_1_subtile_0__pin_O1_7_,
                 top_width_0_height_1_subtile_0__pin_O1_8_,
                 top_width_0_height_1_subtile_0__pin_O1_9_,
                 top_width_0_height_1_subtile_0__pin_O1_10_,
                 top_width_0_height_1_subtile_0__pin_O1_11_,
                 top_width_0_height_2_subtile_0__pin_O2_0_,
                 top_width_0_height_2_subtile_0__pin_O2_1_,
                 top_width_0_height_2_subtile_0__pin_O2_2_,
                 top_width_0_height_2_subtile_0__pin_O2_3_,
                 top_width_0_height_2_subtile_0__pin_O2_4_,
                 top_width_0_height_2_subtile_0__pin_O2_5_,
                 top_width_0_height_2_subtile_0__pin_O2_6_,
                 top_width_0_height_2_subtile_0__pin_O2_7_,
                 top_width_0_height_2_subtile_0__pin_O2_8_,
                 top_width_0_height_2_subtile_0__pin_O2_9_,
                 top_width_0_height_2_subtile_0__pin_O2_10_,
                 top_width_0_height_2_subtile_0__pin_O2_11_,
                 right_width_0_height_0_subtile_0__pin_O0_12_,
                 right_width_0_height_0_subtile_0__pin_O0_13_,
                 right_width_0_height_0_subtile_0__pin_O0_14_,
                 right_width_0_height_0_subtile_0__pin_O0_15_,
                 right_width_0_height_0_subtile_0__pin_O0_16_,
                 right_width_0_height_0_subtile_0__pin_O0_17_,
                 right_width_0_height_0_subtile_0__pin_O0_18_,
                 right_width_0_height_0_subtile_0__pin_O0_19_,
                 right_width_0_height_0_subtile_0__pin_O0_20_,
                 right_width_0_height_0_subtile_0__pin_O0_21_,
                 right_width_0_height_0_subtile_0__pin_O0_22_,
                 right_width_0_height_0_subtile_0__pin_O0_23_,
                 right_width_0_height_0_subtile_0__pin_sc_out_0_,
                 right_width_0_height_0_subtile_0__pin_sc_out_1_,
                 right_width_0_height_0_subtile_0__pin_sc_out_2_,
                 right_width_0_height_0_subtile_0__pin_sc_out_3_,
                 right_width_0_height_0_subtile_0__pin_sc_out_4_,
                 right_width_0_height_0_subtile_0__pin_sc_out_5_,
                 right_width_0_height_1_subtile_0__pin_O1_12_,
                 right_width_0_height_1_subtile_0__pin_O1_13_,
                 right_width_0_height_1_subtile_0__pin_O1_14_,
                 right_width_0_height_1_subtile_0__pin_O1_15_,
                 right_width_0_height_1_subtile_0__pin_O1_16_,
                 right_width_0_height_1_subtile_0__pin_O1_17_,
                 right_width_0_height_1_subtile_0__pin_O1_18_,
                 right_width_0_height_1_subtile_0__pin_O1_19_,
                 right_width_0_height_1_subtile_0__pin_O1_20_,
                 right_width_0_height_1_subtile_0__pin_O1_21_,
                 right_width_0_height_1_subtile_0__pin_O1_22_,
                 right_width_0_height_1_subtile_0__pin_O1_23_,
                 right_width_0_height_2_subtile_0__pin_O2_12_,
                 right_width_0_height_2_subtile_0__pin_O2_13_,
                 right_width_0_height_2_subtile_0__pin_O2_14_,
                 right_width_0_height_2_subtile_0__pin_O2_15_,
                 right_width_0_height_2_subtile_0__pin_O2_16_,
                 right_width_0_height_2_subtile_0__pin_O2_17_,
                 right_width_0_height_2_subtile_0__pin_O2_18_,
                 right_width_0_height_2_subtile_0__pin_O2_19_,
                 right_width_0_height_2_subtile_0__pin_O2_20_,
                 right_width_0_height_2_subtile_0__pin_O2_21_,
                 right_width_0_height_2_subtile_0__pin_O2_22_,
                 right_width_0_height_2_subtile_0__pin_O2_23_,
                 bottom_width_0_height_0_subtile_0__pin_PL_INIT_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ENA_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_REN_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_CLK_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_1_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_1_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_2_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_3_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_4_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_5_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_6_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_7_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_8_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_9_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_10_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_11_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_12_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_13_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_14_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_15_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_16_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_17_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_18_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_19_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_20_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_21_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_22_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_23_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_24_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_25_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_26_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_27_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_28_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_29_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_30_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_31_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_1_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_2_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_3_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_4_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_5_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_6_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_7_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_8_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_9_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_10_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_11_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_12_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_13_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_14_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_15_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_16_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_17_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_18_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_19_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_20_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_21_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_22_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_23_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_24_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_25_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_26_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_27_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_28_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_29_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_30_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_31_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_32_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_33_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_34_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_35_,
                 left_width_0_height_0_subtile_0__pin_sr_out_0_,
                 left_width_0_height_0_subtile_0__pin_sr_out_1_,
                 left_width_0_height_0_subtile_0__pin_sr_out_2_,
                 left_width_0_height_0_subtile_0__pin_sr_out_3_,
                 left_width_0_height_0_subtile_0__pin_sr_out_4_,
                 left_width_0_height_0_subtile_0__pin_sr_out_5_,
                 left_width_0_height_0_subtile_0__pin_plr_o_0_,
                 left_width_0_height_0_subtile_0__pin_plr_o_1_,
                 left_width_0_height_0_subtile_0__pin_plr_o_2_,
                 left_width_0_height_0_subtile_0__pin_plr_o_3_,
                 left_width_0_height_0_subtile_0__pin_plr_o_4_,
                 left_width_0_height_0_subtile_0__pin_plr_o_5_,
                 left_width_0_height_0_subtile_0__pin_plr_o_6_,
                 left_width_0_height_0_subtile_0__pin_plr_o_7_,
                 left_width_0_height_0_subtile_0__pin_plr_o_8_,
                 left_width_0_height_0_subtile_0__pin_plr_o_9_,
                 left_width_0_height_0_subtile_0__pin_plr_o_10_,
                 left_width_0_height_0_subtile_0__pin_plr_o_11_,
                 left_width_0_height_0_subtile_0__pin_plr_o_12_,
                 left_width_0_height_0_subtile_0__pin_plr_o_13_,
                 left_width_0_height_0_subtile_0__pin_plr_o_14_,
                 left_width_0_height_0_subtile_0__pin_plr_o_15_,
                 left_width_0_height_0_subtile_0__pin_plr_o_16_,
                 left_width_0_height_0_subtile_0__pin_plr_o_17_,
                 left_width_0_height_0_subtile_0__pin_plr_o_18_,
                 left_width_0_height_0_subtile_0__pin_plr_o_19_,
                 left_width_0_height_0_subtile_0__pin_plr_o_20_,
                 left_width_0_height_0_subtile_0__pin_plr_o_21_,
                 left_width_0_height_0_subtile_0__pin_plr_o_22_,
                 left_width_0_height_0_subtile_0__pin_plr_o_23_,
                 left_width_0_height_0_subtile_0__pin_plr_o_24_,
                 left_width_0_height_0_subtile_0__pin_plr_o_25_,
                 left_width_0_height_0_subtile_0__pin_plr_o_26_,
                 left_width_0_height_0_subtile_0__pin_plr_o_27_,
                 left_width_0_height_0_subtile_0__pin_plr_o_28_,
                 left_width_0_height_0_subtile_0__pin_plr_o_29_,
                 left_width_0_height_0_subtile_0__pin_plr_o_30_,
                 left_width_0_height_0_subtile_0__pin_plr_o_31_,
                 left_width_0_height_0_subtile_0__pin_plr_o_32_,
                 left_width_0_height_0_subtile_0__pin_plr_o_33_,
                 left_width_0_height_0_subtile_0__pin_plr_o_34_,
                 left_width_0_height_0_subtile_0__pin_plr_o_35_);
//----- GLOBAL PORTS -----
input [0:0] global_resetn;
//----- GLOBAL PORTS -----
input [0:0] scan_en;
//----- GLOBAL PORTS -----
input [0:0] scan_mode;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_INIT_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ENA_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_REN_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_WEN_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_WEN_i_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_12_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_13_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_14_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_15_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_16_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_17_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_18_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_19_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_20_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_21_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_22_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_23_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_24_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_25_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_26_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_27_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_28_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_29_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_30_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_ADDR_i_31_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_12_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_13_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_14_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_15_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_16_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_17_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_18_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_19_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_20_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_21_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_22_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_23_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_24_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_25_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_26_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_27_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_28_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_29_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_30_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_31_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_32_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_33_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_34_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_i_35_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_CLK_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_sr_in_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_sr_in_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_sr_in_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_sr_in_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_sr_in_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_sr_in_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_14_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_15_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_16_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_17_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_18_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_19_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_20_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_21_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_22_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_23_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_24_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_25_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_26_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_27_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_28_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_29_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_30_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_31_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_32_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_33_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_34_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_plr_i_35_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_16_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_17_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_19_;
//----- INPUT PORTS -----
input [0:28] bl;
//----- INPUT PORTS -----
input [0:28] wl;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_23_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_INIT_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ENA_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_REN_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_CLK_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_3_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_5_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_6_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_7_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_8_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_9_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_10_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_11_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_13_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_14_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_15_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_17_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_18_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_19_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_20_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_21_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_22_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_23_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_24_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_25_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_26_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_27_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_28_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_29_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_30_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_31_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_3_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_5_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_6_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_7_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_8_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_9_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_10_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_11_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_13_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_14_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_15_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_17_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_18_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_19_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_20_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_21_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_22_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_23_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_24_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_25_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_26_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_27_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_28_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_29_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_30_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_31_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_32_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_33_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_34_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_35_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_sr_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_sr_out_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_sr_out_2_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_sr_out_3_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_sr_out_4_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_sr_out_5_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_2_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_3_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_4_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_5_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_6_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_7_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_8_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_9_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_10_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_11_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_12_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_13_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_14_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_15_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_16_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_17_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_18_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_19_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_20_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_21_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_22_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_23_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_24_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_25_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_26_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_27_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_28_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_29_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_30_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_31_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_32_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_33_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_34_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_plr_o_35_;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_bram_mode_bram_ logical_tile_bram_mode_bram__0 (
		.global_resetn(global_resetn),
		.scan_en(scan_en),
		.scan_mode(scan_mode),
		.bram_I00({top_width_0_height_0_subtile_0__pin_I00_0_, top_width_0_height_0_subtile_0__pin_I00_1_, top_width_0_height_0_subtile_0__pin_I00_2_, top_width_0_height_0_subtile_0__pin_I00_3_, top_width_0_height_0_subtile_0__pin_I00_4_, top_width_0_height_0_subtile_0__pin_I00_5_, top_width_0_height_0_subtile_0__pin_I00_6_, top_width_0_height_0_subtile_0__pin_I00_7_, top_width_0_height_0_subtile_0__pin_I00_8_, top_width_0_height_0_subtile_0__pin_I00_9_, top_width_0_height_0_subtile_0__pin_I00_10_, top_width_0_height_0_subtile_0__pin_I00_11_}),
		.bram_I10({top_width_0_height_0_subtile_0__pin_I10_0_, top_width_0_height_0_subtile_0__pin_I10_1_, top_width_0_height_0_subtile_0__pin_I10_2_, top_width_0_height_0_subtile_0__pin_I10_3_, top_width_0_height_0_subtile_0__pin_I10_4_, top_width_0_height_0_subtile_0__pin_I10_5_, top_width_0_height_0_subtile_0__pin_I10_6_, top_width_0_height_0_subtile_0__pin_I10_7_, top_width_0_height_0_subtile_0__pin_I10_8_, top_width_0_height_0_subtile_0__pin_I10_9_, top_width_0_height_0_subtile_0__pin_I10_10_, top_width_0_height_0_subtile_0__pin_I10_11_}),
		.bram_I20({right_width_0_height_0_subtile_0__pin_I20_0_, right_width_0_height_0_subtile_0__pin_I20_1_, right_width_0_height_0_subtile_0__pin_I20_2_, right_width_0_height_0_subtile_0__pin_I20_3_, right_width_0_height_0_subtile_0__pin_I20_4_, right_width_0_height_0_subtile_0__pin_I20_5_, right_width_0_height_0_subtile_0__pin_I20_6_, right_width_0_height_0_subtile_0__pin_I20_7_, right_width_0_height_0_subtile_0__pin_I20_8_, right_width_0_height_0_subtile_0__pin_I20_9_, right_width_0_height_0_subtile_0__pin_I20_10_, right_width_0_height_0_subtile_0__pin_I20_11_}),
		.bram_I30({right_width_0_height_0_subtile_0__pin_I30_0_, right_width_0_height_0_subtile_0__pin_I30_1_, right_width_0_height_0_subtile_0__pin_I30_2_, right_width_0_height_0_subtile_0__pin_I30_3_, right_width_0_height_0_subtile_0__pin_I30_4_, right_width_0_height_0_subtile_0__pin_I30_5_, right_width_0_height_0_subtile_0__pin_I30_6_, right_width_0_height_0_subtile_0__pin_I30_7_, right_width_0_height_0_subtile_0__pin_I30_8_, right_width_0_height_0_subtile_0__pin_I30_9_, right_width_0_height_0_subtile_0__pin_I30_10_, right_width_0_height_0_subtile_0__pin_I30_11_}),
		.bram_IS0({top_width_0_height_0_subtile_0__pin_IS0_0_, top_width_0_height_0_subtile_0__pin_IS0_1_, top_width_0_height_0_subtile_0__pin_IS0_2_, right_width_0_height_0_subtile_0__pin_IS0_3_, right_width_0_height_0_subtile_0__pin_IS0_4_, right_width_0_height_0_subtile_0__pin_IS0_5_}),
		.bram_I01({top_width_0_height_1_subtile_0__pin_I01_0_, top_width_0_height_1_subtile_0__pin_I01_1_, top_width_0_height_1_subtile_0__pin_I01_2_, top_width_0_height_1_subtile_0__pin_I01_3_, top_width_0_height_1_subtile_0__pin_I01_4_, top_width_0_height_1_subtile_0__pin_I01_5_, top_width_0_height_1_subtile_0__pin_I01_6_, top_width_0_height_1_subtile_0__pin_I01_7_, top_width_0_height_1_subtile_0__pin_I01_8_, top_width_0_height_1_subtile_0__pin_I01_9_, top_width_0_height_1_subtile_0__pin_I01_10_, top_width_0_height_1_subtile_0__pin_I01_11_}),
		.bram_I11({top_width_0_height_1_subtile_0__pin_I11_0_, top_width_0_height_1_subtile_0__pin_I11_1_, top_width_0_height_1_subtile_0__pin_I11_2_, top_width_0_height_1_subtile_0__pin_I11_3_, top_width_0_height_1_subtile_0__pin_I11_4_, top_width_0_height_1_subtile_0__pin_I11_5_, top_width_0_height_1_subtile_0__pin_I11_6_, top_width_0_height_1_subtile_0__pin_I11_7_, top_width_0_height_1_subtile_0__pin_I11_8_, top_width_0_height_1_subtile_0__pin_I11_9_, top_width_0_height_1_subtile_0__pin_I11_10_, top_width_0_height_1_subtile_0__pin_I11_11_}),
		.bram_I21({right_width_0_height_1_subtile_0__pin_I21_0_, right_width_0_height_1_subtile_0__pin_I21_1_, right_width_0_height_1_subtile_0__pin_I21_2_, right_width_0_height_1_subtile_0__pin_I21_3_, right_width_0_height_1_subtile_0__pin_I21_4_, right_width_0_height_1_subtile_0__pin_I21_5_, right_width_0_height_1_subtile_0__pin_I21_6_, right_width_0_height_1_subtile_0__pin_I21_7_, right_width_0_height_1_subtile_0__pin_I21_8_, right_width_0_height_1_subtile_0__pin_I21_9_, right_width_0_height_1_subtile_0__pin_I21_10_, right_width_0_height_1_subtile_0__pin_I21_11_}),
		.bram_I31({right_width_0_height_1_subtile_0__pin_I31_0_, right_width_0_height_1_subtile_0__pin_I31_1_, right_width_0_height_1_subtile_0__pin_I31_2_, right_width_0_height_1_subtile_0__pin_I31_3_, right_width_0_height_1_subtile_0__pin_I31_4_, right_width_0_height_1_subtile_0__pin_I31_5_, right_width_0_height_1_subtile_0__pin_I31_6_, right_width_0_height_1_subtile_0__pin_I31_7_, right_width_0_height_1_subtile_0__pin_I31_8_, right_width_0_height_1_subtile_0__pin_I31_9_, right_width_0_height_1_subtile_0__pin_I31_10_, right_width_0_height_1_subtile_0__pin_I31_11_}),
		.bram_IS1({top_width_0_height_1_subtile_0__pin_IS1_0_, top_width_0_height_1_subtile_0__pin_IS1_1_, top_width_0_height_1_subtile_0__pin_IS1_2_, right_width_0_height_1_subtile_0__pin_IS1_3_, right_width_0_height_1_subtile_0__pin_IS1_4_, right_width_0_height_1_subtile_0__pin_IS1_5_}),
		.bram_I02({top_width_0_height_2_subtile_0__pin_I02_0_, top_width_0_height_2_subtile_0__pin_I02_1_, top_width_0_height_2_subtile_0__pin_I02_2_, top_width_0_height_2_subtile_0__pin_I02_3_, top_width_0_height_2_subtile_0__pin_I02_4_, top_width_0_height_2_subtile_0__pin_I02_5_, top_width_0_height_2_subtile_0__pin_I02_6_, top_width_0_height_2_subtile_0__pin_I02_7_, top_width_0_height_2_subtile_0__pin_I02_8_, top_width_0_height_2_subtile_0__pin_I02_9_, top_width_0_height_2_subtile_0__pin_I02_10_, top_width_0_height_2_subtile_0__pin_I02_11_}),
		.bram_I12({top_width_0_height_2_subtile_0__pin_I12_0_, top_width_0_height_2_subtile_0__pin_I12_1_, top_width_0_height_2_subtile_0__pin_I12_2_, top_width_0_height_2_subtile_0__pin_I12_3_, top_width_0_height_2_subtile_0__pin_I12_4_, top_width_0_height_2_subtile_0__pin_I12_5_, top_width_0_height_2_subtile_0__pin_I12_6_, top_width_0_height_2_subtile_0__pin_I12_7_, top_width_0_height_2_subtile_0__pin_I12_8_, top_width_0_height_2_subtile_0__pin_I12_9_, top_width_0_height_2_subtile_0__pin_I12_10_, top_width_0_height_2_subtile_0__pin_I12_11_}),
		.bram_I22({right_width_0_height_2_subtile_0__pin_I22_0_, right_width_0_height_2_subtile_0__pin_I22_1_, right_width_0_height_2_subtile_0__pin_I22_2_, right_width_0_height_2_subtile_0__pin_I22_3_, right_width_0_height_2_subtile_0__pin_I22_4_, right_width_0_height_2_subtile_0__pin_I22_5_, right_width_0_height_2_subtile_0__pin_I22_6_, right_width_0_height_2_subtile_0__pin_I22_7_, right_width_0_height_2_subtile_0__pin_I22_8_, right_width_0_height_2_subtile_0__pin_I22_9_, right_width_0_height_2_subtile_0__pin_I22_10_, right_width_0_height_2_subtile_0__pin_I22_11_}),
		.bram_I32({right_width_0_height_2_subtile_0__pin_I32_0_, right_width_0_height_2_subtile_0__pin_I32_1_, right_width_0_height_2_subtile_0__pin_I32_2_, right_width_0_height_2_subtile_0__pin_I32_3_, right_width_0_height_2_subtile_0__pin_I32_4_, right_width_0_height_2_subtile_0__pin_I32_5_, right_width_0_height_2_subtile_0__pin_I32_6_, right_width_0_height_2_subtile_0__pin_I32_7_, right_width_0_height_2_subtile_0__pin_I32_8_, right_width_0_height_2_subtile_0__pin_I32_9_, right_width_0_height_2_subtile_0__pin_I32_10_, right_width_0_height_2_subtile_0__pin_I32_11_}),
		.bram_IS2({top_width_0_height_2_subtile_0__pin_IS2_0_, top_width_0_height_2_subtile_0__pin_IS2_1_, top_width_0_height_2_subtile_0__pin_IS2_2_, right_width_0_height_2_subtile_0__pin_IS2_3_, right_width_0_height_2_subtile_0__pin_IS2_4_, right_width_0_height_2_subtile_0__pin_IS2_5_}),
		.bram_RAM_ID_i({left_width_0_height_1_subtile_0__pin_RAM_ID_i_0_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_1_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_2_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_3_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_4_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_5_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_6_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_7_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_8_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_9_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_10_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_11_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_12_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_13_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_14_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_15_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_16_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_17_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_18_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_19_}),
		.bram_PL_INIT_i(top_width_0_height_2_subtile_0__pin_PL_INIT_i_0_),
		.bram_PL_ENA_i(top_width_0_height_2_subtile_0__pin_PL_ENA_i_0_),
		.bram_PL_REN_i(top_width_0_height_2_subtile_0__pin_PL_REN_i_0_),
		.bram_PL_WEN_i({top_width_0_height_2_subtile_0__pin_PL_WEN_i_0_, top_width_0_height_2_subtile_0__pin_PL_WEN_i_1_}),
		.bram_PL_ADDR_i({top_width_0_height_2_subtile_0__pin_PL_ADDR_i_0_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_1_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_2_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_3_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_4_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_5_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_6_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_7_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_8_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_9_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_10_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_11_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_12_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_13_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_14_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_15_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_16_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_17_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_18_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_19_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_20_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_21_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_22_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_23_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_24_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_25_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_26_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_27_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_28_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_29_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_30_, top_width_0_height_2_subtile_0__pin_PL_ADDR_i_31_}),
		.bram_PL_DATA_i({top_width_0_height_2_subtile_0__pin_PL_DATA_i_0_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_1_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_2_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_3_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_4_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_5_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_6_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_7_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_8_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_9_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_10_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_11_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_12_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_13_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_14_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_15_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_16_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_17_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_18_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_19_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_20_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_21_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_22_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_23_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_24_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_25_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_26_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_27_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_28_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_29_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_30_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_31_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_32_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_33_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_34_, top_width_0_height_2_subtile_0__pin_PL_DATA_i_35_}),
		.bram_sc_in({left_width_0_height_0_subtile_0__pin_sc_in_0_, left_width_0_height_0_subtile_0__pin_sc_in_1_, left_width_0_height_0_subtile_0__pin_sc_in_2_, left_width_0_height_0_subtile_0__pin_sc_in_3_, left_width_0_height_0_subtile_0__pin_sc_in_4_, left_width_0_height_0_subtile_0__pin_sc_in_5_}),
		.bram_sr_in({right_width_0_height_0_subtile_0__pin_sr_in_0_, right_width_0_height_0_subtile_0__pin_sr_in_1_, right_width_0_height_0_subtile_0__pin_sr_in_2_, right_width_0_height_0_subtile_0__pin_sr_in_3_, right_width_0_height_0_subtile_0__pin_sr_in_4_, right_width_0_height_0_subtile_0__pin_sr_in_5_}),
		.bram_plr_i({right_width_0_height_0_subtile_0__pin_plr_i_0_, right_width_0_height_0_subtile_0__pin_plr_i_1_, right_width_0_height_0_subtile_0__pin_plr_i_2_, right_width_0_height_0_subtile_0__pin_plr_i_3_, right_width_0_height_0_subtile_0__pin_plr_i_4_, right_width_0_height_0_subtile_0__pin_plr_i_5_, right_width_0_height_0_subtile_0__pin_plr_i_6_, right_width_0_height_0_subtile_0__pin_plr_i_7_, right_width_0_height_0_subtile_0__pin_plr_i_8_, right_width_0_height_0_subtile_0__pin_plr_i_9_, right_width_0_height_0_subtile_0__pin_plr_i_10_, right_width_0_height_0_subtile_0__pin_plr_i_11_, right_width_0_height_0_subtile_0__pin_plr_i_12_, right_width_0_height_0_subtile_0__pin_plr_i_13_, right_width_0_height_0_subtile_0__pin_plr_i_14_, right_width_0_height_0_subtile_0__pin_plr_i_15_, right_width_0_height_0_subtile_0__pin_plr_i_16_, right_width_0_height_0_subtile_0__pin_plr_i_17_, right_width_0_height_0_subtile_0__pin_plr_i_18_, right_width_0_height_0_subtile_0__pin_plr_i_19_, right_width_0_height_0_subtile_0__pin_plr_i_20_, right_width_0_height_0_subtile_0__pin_plr_i_21_, right_width_0_height_0_subtile_0__pin_plr_i_22_, right_width_0_height_0_subtile_0__pin_plr_i_23_, right_width_0_height_0_subtile_0__pin_plr_i_24_, right_width_0_height_0_subtile_0__pin_plr_i_25_, right_width_0_height_0_subtile_0__pin_plr_i_26_, right_width_0_height_0_subtile_0__pin_plr_i_27_, right_width_0_height_0_subtile_0__pin_plr_i_28_, right_width_0_height_0_subtile_0__pin_plr_i_29_, right_width_0_height_0_subtile_0__pin_plr_i_30_, right_width_0_height_0_subtile_0__pin_plr_i_31_, right_width_0_height_0_subtile_0__pin_plr_i_32_, right_width_0_height_0_subtile_0__pin_plr_i_33_, right_width_0_height_0_subtile_0__pin_plr_i_34_, right_width_0_height_0_subtile_0__pin_plr_i_35_}),
		.bram_PL_CLK_i(top_width_0_height_2_subtile_0__pin_PL_CLK_i_0_),
		.bram_clk({left_width_0_height_0_subtile_0__pin_clk_0_, left_width_0_height_0_subtile_0__pin_clk_1_, left_width_0_height_0_subtile_0__pin_clk_2_, left_width_0_height_0_subtile_0__pin_clk_3_, left_width_0_height_0_subtile_0__pin_clk_4_, left_width_0_height_0_subtile_0__pin_clk_5_, left_width_0_height_0_subtile_0__pin_clk_6_, left_width_0_height_0_subtile_0__pin_clk_7_, left_width_0_height_0_subtile_0__pin_clk_8_, left_width_0_height_0_subtile_0__pin_clk_9_, left_width_0_height_0_subtile_0__pin_clk_10_, left_width_0_height_0_subtile_0__pin_clk_11_, left_width_0_height_0_subtile_0__pin_clk_12_, left_width_0_height_0_subtile_0__pin_clk_13_, left_width_0_height_0_subtile_0__pin_clk_14_, left_width_0_height_0_subtile_0__pin_clk_15_}),
		.bl({bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:28], bl[0:27]}),
		.wl({wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0:1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1:2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2:3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3:4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4:5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5:6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6:7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7:8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8:9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9:10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10:11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11:12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12:13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13:14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14], wl[14:15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15], wl[15:16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16], wl[16:17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17], wl[17:18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18], wl[18:19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19], wl[19:20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20], wl[20:21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21], wl[21:22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22], wl[22:23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23], wl[23:24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24], wl[24:25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25], wl[25:26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26], wl[26:27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27], wl[27:28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28], wl[28]}),
		.bram_O0({top_width_0_height_0_subtile_0__pin_O0_0_, top_width_0_height_0_subtile_0__pin_O0_1_, top_width_0_height_0_subtile_0__pin_O0_2_, top_width_0_height_0_subtile_0__pin_O0_3_, top_width_0_height_0_subtile_0__pin_O0_4_, top_width_0_height_0_subtile_0__pin_O0_5_, top_width_0_height_0_subtile_0__pin_O0_6_, top_width_0_height_0_subtile_0__pin_O0_7_, top_width_0_height_0_subtile_0__pin_O0_8_, top_width_0_height_0_subtile_0__pin_O0_9_, top_width_0_height_0_subtile_0__pin_O0_10_, top_width_0_height_0_subtile_0__pin_O0_11_, right_width_0_height_0_subtile_0__pin_O0_12_, right_width_0_height_0_subtile_0__pin_O0_13_, right_width_0_height_0_subtile_0__pin_O0_14_, right_width_0_height_0_subtile_0__pin_O0_15_, right_width_0_height_0_subtile_0__pin_O0_16_, right_width_0_height_0_subtile_0__pin_O0_17_, right_width_0_height_0_subtile_0__pin_O0_18_, right_width_0_height_0_subtile_0__pin_O0_19_, right_width_0_height_0_subtile_0__pin_O0_20_, right_width_0_height_0_subtile_0__pin_O0_21_, right_width_0_height_0_subtile_0__pin_O0_22_, right_width_0_height_0_subtile_0__pin_O0_23_}),
		.bram_O1({top_width_0_height_1_subtile_0__pin_O1_0_, top_width_0_height_1_subtile_0__pin_O1_1_, top_width_0_height_1_subtile_0__pin_O1_2_, top_width_0_height_1_subtile_0__pin_O1_3_, top_width_0_height_1_subtile_0__pin_O1_4_, top_width_0_height_1_subtile_0__pin_O1_5_, top_width_0_height_1_subtile_0__pin_O1_6_, top_width_0_height_1_subtile_0__pin_O1_7_, top_width_0_height_1_subtile_0__pin_O1_8_, top_width_0_height_1_subtile_0__pin_O1_9_, top_width_0_height_1_subtile_0__pin_O1_10_, top_width_0_height_1_subtile_0__pin_O1_11_, right_width_0_height_1_subtile_0__pin_O1_12_, right_width_0_height_1_subtile_0__pin_O1_13_, right_width_0_height_1_subtile_0__pin_O1_14_, right_width_0_height_1_subtile_0__pin_O1_15_, right_width_0_height_1_subtile_0__pin_O1_16_, right_width_0_height_1_subtile_0__pin_O1_17_, right_width_0_height_1_subtile_0__pin_O1_18_, right_width_0_height_1_subtile_0__pin_O1_19_, right_width_0_height_1_subtile_0__pin_O1_20_, right_width_0_height_1_subtile_0__pin_O1_21_, right_width_0_height_1_subtile_0__pin_O1_22_, right_width_0_height_1_subtile_0__pin_O1_23_}),
		.bram_O2({top_width_0_height_2_subtile_0__pin_O2_0_, top_width_0_height_2_subtile_0__pin_O2_1_, top_width_0_height_2_subtile_0__pin_O2_2_, top_width_0_height_2_subtile_0__pin_O2_3_, top_width_0_height_2_subtile_0__pin_O2_4_, top_width_0_height_2_subtile_0__pin_O2_5_, top_width_0_height_2_subtile_0__pin_O2_6_, top_width_0_height_2_subtile_0__pin_O2_7_, top_width_0_height_2_subtile_0__pin_O2_8_, top_width_0_height_2_subtile_0__pin_O2_9_, top_width_0_height_2_subtile_0__pin_O2_10_, top_width_0_height_2_subtile_0__pin_O2_11_, right_width_0_height_2_subtile_0__pin_O2_12_, right_width_0_height_2_subtile_0__pin_O2_13_, right_width_0_height_2_subtile_0__pin_O2_14_, right_width_0_height_2_subtile_0__pin_O2_15_, right_width_0_height_2_subtile_0__pin_O2_16_, right_width_0_height_2_subtile_0__pin_O2_17_, right_width_0_height_2_subtile_0__pin_O2_18_, right_width_0_height_2_subtile_0__pin_O2_19_, right_width_0_height_2_subtile_0__pin_O2_20_, right_width_0_height_2_subtile_0__pin_O2_21_, right_width_0_height_2_subtile_0__pin_O2_22_, right_width_0_height_2_subtile_0__pin_O2_23_}),
		.bram_PL_INIT_o(bottom_width_0_height_0_subtile_0__pin_PL_INIT_o_0_),
		.bram_PL_ENA_o(bottom_width_0_height_0_subtile_0__pin_PL_ENA_o_0_),
		.bram_PL_REN_o(bottom_width_0_height_0_subtile_0__pin_PL_REN_o_0_),
		.bram_PL_CLK_o(bottom_width_0_height_0_subtile_0__pin_PL_CLK_o_0_),
		.bram_PL_WEN_o({bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_0_, bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_1_}),
		.bram_PL_ADDR_o({bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_0_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_1_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_2_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_3_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_4_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_5_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_6_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_7_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_8_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_9_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_10_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_11_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_12_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_13_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_14_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_15_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_16_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_17_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_18_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_19_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_20_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_21_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_22_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_23_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_24_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_25_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_26_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_27_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_28_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_29_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_30_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_31_}),
		.bram_PL_DATA_o({bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_0_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_1_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_2_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_3_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_4_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_5_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_6_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_7_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_8_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_9_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_10_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_11_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_12_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_13_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_14_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_15_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_16_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_17_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_18_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_19_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_20_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_21_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_22_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_23_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_24_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_25_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_26_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_27_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_28_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_29_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_30_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_31_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_32_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_33_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_34_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_35_}),
		.bram_sc_out({right_width_0_height_0_subtile_0__pin_sc_out_0_, right_width_0_height_0_subtile_0__pin_sc_out_1_, right_width_0_height_0_subtile_0__pin_sc_out_2_, right_width_0_height_0_subtile_0__pin_sc_out_3_, right_width_0_height_0_subtile_0__pin_sc_out_4_, right_width_0_height_0_subtile_0__pin_sc_out_5_}),
		.bram_sr_out({left_width_0_height_0_subtile_0__pin_sr_out_0_, left_width_0_height_0_subtile_0__pin_sr_out_1_, left_width_0_height_0_subtile_0__pin_sr_out_2_, left_width_0_height_0_subtile_0__pin_sr_out_3_, left_width_0_height_0_subtile_0__pin_sr_out_4_, left_width_0_height_0_subtile_0__pin_sr_out_5_}),
		.bram_plr_o({left_width_0_height_0_subtile_0__pin_plr_o_0_, left_width_0_height_0_subtile_0__pin_plr_o_1_, left_width_0_height_0_subtile_0__pin_plr_o_2_, left_width_0_height_0_subtile_0__pin_plr_o_3_, left_width_0_height_0_subtile_0__pin_plr_o_4_, left_width_0_height_0_subtile_0__pin_plr_o_5_, left_width_0_height_0_subtile_0__pin_plr_o_6_, left_width_0_height_0_subtile_0__pin_plr_o_7_, left_width_0_height_0_subtile_0__pin_plr_o_8_, left_width_0_height_0_subtile_0__pin_plr_o_9_, left_width_0_height_0_subtile_0__pin_plr_o_10_, left_width_0_height_0_subtile_0__pin_plr_o_11_, left_width_0_height_0_subtile_0__pin_plr_o_12_, left_width_0_height_0_subtile_0__pin_plr_o_13_, left_width_0_height_0_subtile_0__pin_plr_o_14_, left_width_0_height_0_subtile_0__pin_plr_o_15_, left_width_0_height_0_subtile_0__pin_plr_o_16_, left_width_0_height_0_subtile_0__pin_plr_o_17_, left_width_0_height_0_subtile_0__pin_plr_o_18_, left_width_0_height_0_subtile_0__pin_plr_o_19_, left_width_0_height_0_subtile_0__pin_plr_o_20_, left_width_0_height_0_subtile_0__pin_plr_o_21_, left_width_0_height_0_subtile_0__pin_plr_o_22_, left_width_0_height_0_subtile_0__pin_plr_o_23_, left_width_0_height_0_subtile_0__pin_plr_o_24_, left_width_0_height_0_subtile_0__pin_plr_o_25_, left_width_0_height_0_subtile_0__pin_plr_o_26_, left_width_0_height_0_subtile_0__pin_plr_o_27_, left_width_0_height_0_subtile_0__pin_plr_o_28_, left_width_0_height_0_subtile_0__pin_plr_o_29_, left_width_0_height_0_subtile_0__pin_plr_o_30_, left_width_0_height_0_subtile_0__pin_plr_o_31_, left_width_0_height_0_subtile_0__pin_plr_o_32_, left_width_0_height_0_subtile_0__pin_plr_o_33_, left_width_0_height_0_subtile_0__pin_plr_o_34_, left_width_0_height_0_subtile_0__pin_plr_o_35_}));

endmodule
// ----- END Verilog module for grid_bram -----

//----- Default net type -----
`default_nettype none



// ----- END Grid Verilog module: grid_bram -----

