//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[10][8]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_10__8_ -----
module sb_10__8_(chany_bottom_in,
                 bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_,
                 chanx_left_in,
                 left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_,
                 bl,
                 wl,
                 chany_bottom_out,
                 chanx_left_out);
//----- INPUT PORTS -----
input [0:79] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:79] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:19] bl;
//----- INPUT PORTS -----
input [0:18] wl;
//----- OUTPUT PORTS -----
output [0:79] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:79] chanx_left_out;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_L1SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_10_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_11_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_6_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_7_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_8_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_9_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_30_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_31_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_14_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_15_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_16_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_17_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_17_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_18_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_18_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_19_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_19_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_20_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_20_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_21_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_21_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_22_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_22_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_23_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_23_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_24_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_24_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_25_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_25_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_26_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_26_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_27_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_27_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_28_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_28_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_29_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_29_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_30_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_30_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_31_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_31_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_16_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_16_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_17_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_17_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_18_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_18_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_19_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_19_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_20_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_20_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_21_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_21_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_22_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_22_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_23_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_23_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_24_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_24_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_25_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_25_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_26_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_26_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_27_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_27_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_28_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_28_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_29_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_29_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_30_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_30_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_31_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_31_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[12] = chany_bottom_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[15] = chany_bottom_in[14];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_1 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, chanx_left_in[1]}),
		.sram(mux_tree_tapbuf_L1SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_3 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, chanx_left_in[2]}),
		.sram(mux_tree_tapbuf_L1SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_5 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, chanx_left_in[3]}),
		.sram(mux_tree_tapbuf_L1SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_2_sram_inv[0:2]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_7 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, chanx_left_in[4]}),
		.sram(mux_tree_tapbuf_L1SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_3_sram_inv[0:2]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_9 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[5]}),
		.sram(mux_tree_tapbuf_L1SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_4_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_11 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[6]}),
		.sram(mux_tree_tapbuf_L1SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_5_sram_inv[0:2]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_13 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[7]}),
		.sram(mux_tree_tapbuf_L1SB_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_6_sram_inv[0:2]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_15 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[8]}),
		.sram(mux_tree_tapbuf_L1SB_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_7_sram_inv[0:2]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_17 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[9]}),
		.sram(mux_tree_tapbuf_L1SB_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_8_sram_inv[0:2]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_19 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[10]}),
		.sram(mux_tree_tapbuf_L1SB_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_9_sram_inv[0:2]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_21 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[11]}),
		.sram(mux_tree_tapbuf_L1SB_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_10_sram_inv[0:2]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_23 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[12]}),
		.sram(mux_tree_tapbuf_L1SB_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_11_sram_inv[0:2]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_1 (
		.bl(bl[0:2]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_3 (
		.bl(bl[3:5]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_5 (
		.bl(bl[6:8]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_7 (
		.bl(bl[9:11]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_9 (
		.bl(bl[12:14]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_11 (
		.bl(bl[15:17]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_13 (
		.bl({bl[18:19], bl[0]}),
		.wl({wl[0], wl[0:1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_15 (
		.bl(bl[1:3]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_17 (
		.bl(bl[4:6]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_19 (
		.bl(bl[7:9]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_21 (
		.bl(bl[10:12]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_23 (
		.bl(bl[13:15]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size4 mux_bottom_track_25 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, chanx_left_in[13]}),
		.sram(mux_tree_tapbuf_L1SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_0_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_L1SB_size4 mux_bottom_track_27 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, chanx_left_in[14]}),
		.sram(mux_tree_tapbuf_L1SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_1_sram_inv[0:1]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_L1SB_size4 mux_bottom_track_29 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, chanx_left_in[15]}),
		.sram(mux_tree_tapbuf_L1SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_2_sram_inv[0:1]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_L1SB_size4 mux_bottom_track_31 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, chanx_left_in[16]}),
		.sram(mux_tree_tapbuf_L1SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_3_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_L1SB_size4_mem mem_bottom_track_25 (
		.bl(bl[16:17]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_bottom_track_27 (
		.bl(bl[18:19]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_bottom_track_29 (
		.bl(bl[0:1]),
		.wl({wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_bottom_track_31 (
		.bl(bl[2:3]),
		.wl({wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_33 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[17]}),
		.sram(mux_tree_tapbuf_L4SB_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_0_sram_inv[0:3]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_35 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[18]}),
		.sram(mux_tree_tapbuf_L4SB_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_1_sram_inv[0:3]),
		.out(chany_bottom_out[17]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_37 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[19]}),
		.sram(mux_tree_tapbuf_L4SB_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_2_sram_inv[0:3]),
		.out(chany_bottom_out[18]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_39 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[20]}),
		.sram(mux_tree_tapbuf_L4SB_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_3_sram_inv[0:3]),
		.out(chany_bottom_out[19]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_49 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[25]}),
		.sram(mux_tree_tapbuf_L4SB_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_4_sram_inv[0:3]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_51 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[26]}),
		.sram(mux_tree_tapbuf_L4SB_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_5_sram_inv[0:3]),
		.out(chany_bottom_out[25]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_53 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[27]}),
		.sram(mux_tree_tapbuf_L4SB_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_6_sram_inv[0:3]),
		.out(chany_bottom_out[26]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_55 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[28]}),
		.sram(mux_tree_tapbuf_L4SB_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_7_sram_inv[0:3]),
		.out(chany_bottom_out[27]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_65 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[33]}),
		.sram(mux_tree_tapbuf_L4SB_size9_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_8_sram_inv[0:3]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_67 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[34]}),
		.sram(mux_tree_tapbuf_L4SB_size9_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_9_sram_inv[0:3]),
		.out(chany_bottom_out[33]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_69 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[35]}),
		.sram(mux_tree_tapbuf_L4SB_size9_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_10_sram_inv[0:3]),
		.out(chany_bottom_out[34]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_71 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[36]}),
		.sram(mux_tree_tapbuf_L4SB_size9_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_11_sram_inv[0:3]),
		.out(chany_bottom_out[35]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_81 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size9_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_12_sram_inv[0:3]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_83 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size9_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_13_sram_inv[0:3]),
		.out(chany_bottom_out[41]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_85 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_L4SB_size9_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_14_sram_inv[0:3]),
		.out(chany_bottom_out[42]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_87 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size9_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_15_sram_inv[0:3]),
		.out(chany_bottom_out[43]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_97 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size9_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_16_sram_inv[0:3]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_99 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size9_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_17_sram_inv[0:3]),
		.out(chany_bottom_out[49]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_101 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size9_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_18_sram_inv[0:3]),
		.out(chany_bottom_out[50]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_103 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size9_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_19_sram_inv[0:3]),
		.out(chany_bottom_out[51]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_113 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size9_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_20_sram_inv[0:3]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_115 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L4SB_size9_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_21_sram_inv[0:3]),
		.out(chany_bottom_out[57]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_117 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size9_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_22_sram_inv[0:3]),
		.out(chany_bottom_out[58]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_119 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size9_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_23_sram_inv[0:3]),
		.out(chany_bottom_out[59]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_129 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size9_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_24_sram_inv[0:3]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_131 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L4SB_size9_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_25_sram_inv[0:3]),
		.out(chany_bottom_out[65]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_133 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size9_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_26_sram_inv[0:3]),
		.out(chany_bottom_out[66]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_135 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size9_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_27_sram_inv[0:3]),
		.out(chany_bottom_out[67]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_145 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size9_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_28_sram_inv[0:3]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_147 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L4SB_size9_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_29_sram_inv[0:3]),
		.out(chany_bottom_out[73]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_149 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size9_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_30_sram_inv[0:3]),
		.out(chany_bottom_out[74]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_151 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L4SB_size9_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_31_sram_inv[0:3]),
		.out(chany_bottom_out[75]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_33 (
		.bl(bl[4:7]),
		.wl({wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_35 (
		.bl(bl[8:11]),
		.wl({wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_37 (
		.bl(bl[12:15]),
		.wl({wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_39 (
		.bl(bl[16:19]),
		.wl({wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_49 (
		.bl(bl[12:15]),
		.wl({wl[3], wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_51 (
		.bl(bl[16:19]),
		.wl({wl[3], wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_53 (
		.bl(bl[0:3]),
		.wl({wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_55 (
		.bl(bl[4:7]),
		.wl({wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_65 (
		.bl(bl[0:3]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_67 (
		.bl(bl[4:7]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_69 (
		.bl(bl[8:11]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_71 (
		.bl(bl[12:15]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_81 (
		.bl(bl[8:11]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_83 (
		.bl(bl[12:15]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_85 (
		.bl(bl[16:19]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_87 (
		.bl(bl[0:3]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_15_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_97 (
		.bl(bl[16:19]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_16_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_99 (
		.bl(bl[0:3]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_17_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_101 (
		.bl(bl[4:7]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_18_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_103 (
		.bl(bl[8:11]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_19_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_113 (
		.bl(bl[4:7]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_20_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_115 (
		.bl(bl[8:11]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_21_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_117 (
		.bl(bl[12:15]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_22_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_119 (
		.bl(bl[16:19]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_23_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_129 (
		.bl(bl[12:15]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_24_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_131 (
		.bl(bl[16:19]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_25_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_133 (
		.bl(bl[0:3]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_26_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_135 (
		.bl(bl[4:7]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_27_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_145 (
		.bl(bl[0:3]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_28_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_147 (
		.bl(bl[4:7]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_29_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_149 (
		.bl(bl[8:11]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_30_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_151 (
		.bl(bl[12:15]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size9_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_31_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_41 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[21]}),
		.sram(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_43 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[22]}),
		.sram(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]),
		.out(chany_bottom_out[21]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_45 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[23]}),
		.sram(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]),
		.out(chany_bottom_out[22]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_47 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[24]}),
		.sram(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]),
		.out(chany_bottom_out[23]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_57 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[29]}),
		.sram(mux_tree_tapbuf_L4SB_size8_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_4_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_59 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[30]}),
		.sram(mux_tree_tapbuf_L4SB_size8_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_5_sram_inv[0:2]),
		.out(chany_bottom_out[29]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_61 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[31]}),
		.sram(mux_tree_tapbuf_L4SB_size8_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_6_sram_inv[0:2]),
		.out(chany_bottom_out[30]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_63 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[32]}),
		.sram(mux_tree_tapbuf_L4SB_size8_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_7_sram_inv[0:2]),
		.out(chany_bottom_out[31]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_73 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size8_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_8_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_75 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size8_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_9_sram_inv[0:2]),
		.out(chany_bottom_out[37]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_77 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[39]}),
		.sram(mux_tree_tapbuf_L4SB_size8_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_10_sram_inv[0:2]),
		.out(chany_bottom_out[38]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_79 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size8_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_11_sram_inv[0:2]),
		.out(chany_bottom_out[39]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_89 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size8_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_12_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_91 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size8_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_13_sram_inv[0:2]),
		.out(chany_bottom_out[45]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_93 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size8_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_14_sram_inv[0:2]),
		.out(chany_bottom_out[46]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_95 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size8_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_15_sram_inv[0:2]),
		.out(chany_bottom_out[47]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_105 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size8_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_16_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_107 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size8_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_17_sram_inv[0:2]),
		.out(chany_bottom_out[53]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_109 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size8_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_18_sram_inv[0:2]),
		.out(chany_bottom_out[54]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_111 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size8_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_19_sram_inv[0:2]),
		.out(chany_bottom_out[55]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_121 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size8_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_20_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_123 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L4SB_size8_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_21_sram_inv[0:2]),
		.out(chany_bottom_out[61]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_125 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size8_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_22_sram_inv[0:2]),
		.out(chany_bottom_out[62]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_127 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size8_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_23_sram_inv[0:2]),
		.out(chany_bottom_out[63]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_137 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size8_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_24_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_139 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L4SB_size8_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_25_sram_inv[0:2]),
		.out(chany_bottom_out[69]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_141 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size8_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_26_sram_inv[0:2]),
		.out(chany_bottom_out[70]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_143 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size8_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_27_sram_inv[0:2]),
		.out(chany_bottom_out[71]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_153 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L4SB_size8_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_28_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_155 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L4SB_size8_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_29_sram_inv[0:2]),
		.out(chany_bottom_out[77]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_157 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size8_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_30_sram_inv[0:2]),
		.out(chany_bottom_out[78]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_159 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[0]}),
		.sram(mux_tree_tapbuf_L4SB_size8_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_31_sram_inv[0:2]),
		.out(chany_bottom_out[79]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_41 (
		.bl(bl[0:2]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_43 (
		.bl(bl[3:5]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_45 (
		.bl(bl[6:8]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_47 (
		.bl(bl[9:11]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_57 (
		.bl(bl[8:10]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_59 (
		.bl(bl[11:13]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_61 (
		.bl(bl[14:16]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_63 (
		.bl(bl[17:19]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_73 (
		.bl(bl[16:18]),
		.wl({wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_75 (
		.bl({bl[19], bl[0:1]}),
		.wl({wl[5:6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_77 (
		.bl(bl[2:4]),
		.wl({wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_79 (
		.bl(bl[5:7]),
		.wl({wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_89 (
		.bl(bl[4:6]),
		.wl({wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_91 (
		.bl(bl[7:9]),
		.wl({wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_93 (
		.bl(bl[10:12]),
		.wl({wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_14_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_95 (
		.bl(bl[13:15]),
		.wl({wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_15_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_105 (
		.bl(bl[12:14]),
		.wl({wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_16_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_107 (
		.bl(bl[15:17]),
		.wl({wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_17_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_109 (
		.bl({bl[18:19], bl[0]}),
		.wl({wl[8], wl[8:9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_18_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_111 (
		.bl(bl[1:3]),
		.wl({wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_19_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_121 (
		.bl(bl[0:2]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_20_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_123 (
		.bl(bl[3:5]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_21_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_125 (
		.bl(bl[6:8]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_22_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_127 (
		.bl(bl[9:11]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_23_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_137 (
		.bl(bl[8:10]),
		.wl({wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_24_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_139 (
		.bl(bl[11:13]),
		.wl({wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_25_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_141 (
		.bl(bl[14:16]),
		.wl({wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_26_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_143 (
		.bl(bl[17:19]),
		.wl({wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_27_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_153 (
		.bl(bl[16:18]),
		.wl({wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_28_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_155 (
		.bl({bl[19], bl[0:1]}),
		.wl({wl[12:13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_29_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_157 (
		.bl(bl[2:4]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_30_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_159 (
		.bl(bl[5:7]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size8_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_31_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_1 (
		.in({chany_bottom_in[79], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_0_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_0_sram_inv),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_3 (
		.in({chany_bottom_in[0], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_1_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_1_sram_inv),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_5 (
		.in({chany_bottom_in[1], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_2_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_2_sram_inv),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_7 (
		.in({chany_bottom_in[2], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_3_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_3_sram_inv),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_9 (
		.in({chany_bottom_in[3], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_4_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_4_sram_inv),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_11 (
		.in({chany_bottom_in[4], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_5_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_5_sram_inv),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_13 (
		.in({chany_bottom_in[5], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_6_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_6_sram_inv),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_15 (
		.in({chany_bottom_in[6], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_7_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_7_sram_inv),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_17 (
		.in({chany_bottom_in[7], left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_8_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_8_sram_inv),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_19 (
		.in({chany_bottom_in[8], left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_9_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_9_sram_inv),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_21 (
		.in({chany_bottom_in[9], left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_10_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_10_sram_inv),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_L1SB_size2 mux_left_track_23 (
		.in({chany_bottom_in[10], left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size2_11_sram),
		.sram_inv(mux_tree_tapbuf_L1SB_size2_11_sram_inv),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_1 (
		.bl(bl[8]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_0_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_0_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_3 (
		.bl(bl[9]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_1_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_1_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_5 (
		.bl(bl[10]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_2_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_2_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_7 (
		.bl(bl[11]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_3_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_3_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_9 (
		.bl(bl[12]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_4_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_4_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_11 (
		.bl(bl[13]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_5_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_5_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_13 (
		.bl(bl[14]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_6_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_6_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_15 (
		.bl(bl[15]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_7_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_7_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_17 (
		.bl(bl[16]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_8_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_8_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_19 (
		.bl(bl[17]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_9_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_9_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_21 (
		.bl(bl[18]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_10_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_10_sram_inv));

	mux_tree_tapbuf_L1SB_size2_mem mem_left_track_23 (
		.bl(bl[19]),
		.wl(wl[13]),
		.mem_out(mux_tree_tapbuf_L1SB_size2_11_sram),
		.mem_outb(mux_tree_tapbuf_L1SB_size2_11_sram_inv));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_33 (
		.in({chany_bottom_in[15], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_35 (
		.in({chany_bottom_in[16], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_37 (
		.in({chany_bottom_in[17], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_39 (
		.in({chany_bottom_in[18], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_49 (
		.in({chany_bottom_in[23], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_51 (
		.in({chany_bottom_in[24], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_53 (
		.in({chany_bottom_in[25], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_55 (
		.in({chany_bottom_in[26], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_65 (
		.in({chany_bottom_in[31], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_67 (
		.in({chany_bottom_in[32], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_69 (
		.in({chany_bottom_in[33], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_71 (
		.in({chany_bottom_in[34], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_81 (
		.in({chany_bottom_in[39], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_83 (
		.in({chany_bottom_in[40], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_85 (
		.in({chany_bottom_in[41], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_87 (
		.in({chany_bottom_in[42], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_97 (
		.in({chany_bottom_in[47], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_99 (
		.in({chany_bottom_in[48], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_101 (
		.in({chany_bottom_in[49], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_103 (
		.in({chany_bottom_in[50], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_113 (
		.in({chany_bottom_in[55], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_115 (
		.in({chany_bottom_in[56], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_117 (
		.in({chany_bottom_in[57], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_119 (
		.in({chany_bottom_in[58], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_129 (
		.in({chany_bottom_in[63], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_131 (
		.in({chany_bottom_in[64], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_133 (
		.in({chany_bottom_in[65], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_135 (
		.in({chany_bottom_in[66], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_145 (
		.in({chany_bottom_in[71], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_147 (
		.in({chany_bottom_in[72], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]),
		.out(chanx_left_out[73]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_149 (
		.in({chany_bottom_in[73], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_30_sram_inv[0:1]),
		.out(chanx_left_out[74]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_151 (
		.in({chany_bottom_in[74], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_31_sram_inv[0:1]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_33 (
		.bl(bl[0:1]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_35 (
		.bl(bl[2:3]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_37 (
		.bl(bl[4:5]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_39 (
		.bl(bl[6:7]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_49 (
		.bl(bl[12:13]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_51 (
		.bl(bl[14:15]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_53 (
		.bl(bl[16:17]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_55 (
		.bl(bl[18:19]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_65 (
		.bl(bl[4:5]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_67 (
		.bl(bl[6:7]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_69 (
		.bl(bl[8:9]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_71 (
		.bl(bl[10:11]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_81 (
		.bl(bl[16:17]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_83 (
		.bl(bl[18:19]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_85 (
		.bl(bl[0:1]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_87 (
		.bl(bl[2:3]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_97 (
		.bl(bl[8:9]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_99 (
		.bl(bl[10:11]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_101 (
		.bl(bl[12:13]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_103 (
		.bl(bl[14:15]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_113 (
		.bl(bl[0:1]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_115 (
		.bl(bl[2:3]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_117 (
		.bl(bl[4:5]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_119 (
		.bl(bl[6:7]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_129 (
		.bl(bl[12:13]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_131 (
		.bl(bl[14:15]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_133 (
		.bl(bl[16:17]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_135 (
		.bl(bl[18:19]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_145 (
		.bl(bl[4:5]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_147 (
		.bl(bl[6:7]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_149 (
		.bl(bl[8:9]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_151 (
		.bl(bl[10:11]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_41 (
		.in({chany_bottom_in[19], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_0_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_0_sram_inv),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_43 (
		.in({chany_bottom_in[20], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_1_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_1_sram_inv),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_45 (
		.in({chany_bottom_in[21], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_2_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_2_sram_inv),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_47 (
		.in({chany_bottom_in[22], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_3_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_3_sram_inv),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_57 (
		.in({chany_bottom_in[27], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_4_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_4_sram_inv),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_59 (
		.in({chany_bottom_in[28], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_5_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_5_sram_inv),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_61 (
		.in({chany_bottom_in[29], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_6_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_6_sram_inv),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_63 (
		.in({chany_bottom_in[30], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_7_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_7_sram_inv),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_73 (
		.in({chany_bottom_in[35], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_8_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_8_sram_inv),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_75 (
		.in({chany_bottom_in[36], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_9_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_9_sram_inv),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_77 (
		.in({chany_bottom_in[37], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_10_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_10_sram_inv),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_79 (
		.in({chany_bottom_in[38], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_11_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_11_sram_inv),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_89 (
		.in({chany_bottom_in[43], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_12_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_12_sram_inv),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_91 (
		.in({chany_bottom_in[44], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_13_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_13_sram_inv),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_93 (
		.in({chany_bottom_in[45], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_14_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_14_sram_inv),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_95 (
		.in({chany_bottom_in[46], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_15_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_15_sram_inv),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_105 (
		.in({chany_bottom_in[51], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_16_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_16_sram_inv),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_107 (
		.in({chany_bottom_in[52], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_17_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_17_sram_inv),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_109 (
		.in({chany_bottom_in[53], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_18_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_18_sram_inv),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_111 (
		.in({chany_bottom_in[54], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_19_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_19_sram_inv),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_121 (
		.in({chany_bottom_in[59], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_20_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_20_sram_inv),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_123 (
		.in({chany_bottom_in[60], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_21_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_21_sram_inv),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_125 (
		.in({chany_bottom_in[61], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_22_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_22_sram_inv),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_127 (
		.in({chany_bottom_in[62], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_23_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_23_sram_inv),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_137 (
		.in({chany_bottom_in[67], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_24_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_24_sram_inv),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_139 (
		.in({chany_bottom_in[68], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_25_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_25_sram_inv),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_141 (
		.in({chany_bottom_in[69], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_26_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_26_sram_inv),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_143 (
		.in({chany_bottom_in[70], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_27_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_27_sram_inv),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_153 (
		.in({chany_bottom_in[75], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_28_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_28_sram_inv),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_155 (
		.in({chany_bottom_in[76], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_29_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_29_sram_inv),
		.out(chanx_left_out[77]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_157 (
		.in({chany_bottom_in[77], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_30_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_30_sram_inv),
		.out(chanx_left_out[78]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_159 (
		.in({chany_bottom_in[78], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_31_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_31_sram_inv),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_41 (
		.bl(bl[8]),
		.wl(wl[14]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_0_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_0_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_43 (
		.bl(bl[9]),
		.wl(wl[14]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_1_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_1_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_45 (
		.bl(bl[10]),
		.wl(wl[14]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_2_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_2_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_47 (
		.bl(bl[11]),
		.wl(wl[14]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_3_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_3_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_57 (
		.bl(bl[0]),
		.wl(wl[15]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_4_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_4_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_59 (
		.bl(bl[1]),
		.wl(wl[15]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_5_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_5_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_61 (
		.bl(bl[2]),
		.wl(wl[15]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_6_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_6_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_63 (
		.bl(bl[3]),
		.wl(wl[15]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_7_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_7_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_73 (
		.bl(bl[12]),
		.wl(wl[15]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_8_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_8_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_75 (
		.bl(bl[13]),
		.wl(wl[15]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_9_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_9_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_77 (
		.bl(bl[14]),
		.wl(wl[15]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_10_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_10_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_79 (
		.bl(bl[15]),
		.wl(wl[15]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_11_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_11_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_89 (
		.bl(bl[4]),
		.wl(wl[16]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_12_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_12_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_91 (
		.bl(bl[5]),
		.wl(wl[16]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_13_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_13_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_93 (
		.bl(bl[6]),
		.wl(wl[16]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_14_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_14_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_95 (
		.bl(bl[7]),
		.wl(wl[16]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_15_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_15_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_105 (
		.bl(bl[16]),
		.wl(wl[16]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_16_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_16_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_107 (
		.bl(bl[17]),
		.wl(wl[16]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_17_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_17_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_109 (
		.bl(bl[18]),
		.wl(wl[16]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_18_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_18_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_111 (
		.bl(bl[19]),
		.wl(wl[16]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_19_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_19_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_121 (
		.bl(bl[8]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_20_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_20_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_123 (
		.bl(bl[9]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_21_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_21_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_125 (
		.bl(bl[10]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_22_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_22_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_127 (
		.bl(bl[11]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_23_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_23_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_137 (
		.bl(bl[0]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_24_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_24_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_139 (
		.bl(bl[1]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_25_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_25_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_141 (
		.bl(bl[2]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_26_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_26_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_143 (
		.bl(bl[3]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_27_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_27_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_153 (
		.bl(bl[12]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_28_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_28_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_155 (
		.bl(bl[13]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_29_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_29_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_157 (
		.bl(bl[14]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_30_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_30_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_159 (
		.bl(bl[15]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_31_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_31_sram_inv));

endmodule
// ----- END Verilog module for sb_10__8_ -----

//----- Default net type -----
`default_nettype none



