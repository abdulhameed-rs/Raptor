//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[10][1]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_10__1_ -----
module sb_10__1_(chany_top_in,
                 top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_,
                 top_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_,
                 chany_bottom_in,
                 bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_,
                 chanx_left_in,
                 left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_,
                 bl,
                 wl,
                 chany_top_out,
                 chany_bottom_out,
                 chanx_left_out);
//----- INPUT PORTS -----
input [0:79] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:79] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:79] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:19] bl;
//----- INPUT PORTS -----
input [0:19] wl;
//----- OUTPUT PORTS -----
output [0:79] chany_top_out;
//----- OUTPUT PORTS -----
output [0:79] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:79] chanx_left_out;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_L1SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size7_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size7_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size7_2_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size7_3_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size7_4_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_10_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_11_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_12_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_13_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_2_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_3_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_4_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_5_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_6_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_7_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_8_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_9_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_0_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_10_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_11_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_12_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_1_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_2_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_3_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_4_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_5_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_6_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_7_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_8_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_9_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_16_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_16_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_17_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_17_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_8_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L1SB_size9 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, chany_bottom_in[16], chany_bottom_in[58], chanx_left_in[0], chanx_left_in[32], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L1SB_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_0_sram_inv[0:3]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_1 (
		.in({chany_top_in[16], chany_top_in[58], bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, chanx_left_in[1], chanx_left_in[33], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L1SB_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_1_sram_inv[0:3]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_3 (
		.in({chany_top_in[17], chany_top_in[60], bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, chanx_left_in[2], chanx_left_in[34], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L1SB_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_2_sram_inv[0:3]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_5 (
		.in({chany_top_in[18], chany_top_in[61], bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, chanx_left_in[3], chanx_left_in[35], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L1SB_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_3_sram_inv[0:3]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_7 (
		.in({chany_top_in[20], chany_top_in[62], bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, chanx_left_in[4], chanx_left_in[36], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L1SB_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_4_sram_inv[0:3]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_9 (
		.in({chany_top_in[21], chany_top_in[64], bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[5], chanx_left_in[37], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L1SB_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_5_sram_inv[0:3]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_11 (
		.in({chany_top_in[22], chany_top_in[65], bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[6], chanx_left_in[38], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L1SB_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_6_sram_inv[0:3]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_13 (
		.in({chany_top_in[24], chany_top_in[66], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[7], chanx_left_in[39], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L1SB_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_7_sram_inv[0:3]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_15 (
		.in({chany_top_in[25], chany_top_in[68], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[8], chanx_left_in[40], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size9_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_8_sram_inv[0:3]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_17 (
		.in({chany_top_in[26], chany_top_in[69], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[9], chanx_left_in[41], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size9_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_9_sram_inv[0:3]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_19 (
		.in({chany_top_in[28], chany_top_in[70], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[10], chanx_left_in[42], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L1SB_size9_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_10_sram_inv[0:3]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_21 (
		.in({chany_top_in[29], chany_top_in[72], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[11], chanx_left_in[43], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L1SB_size9_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_11_sram_inv[0:3]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_23 (
		.in({chany_top_in[30], chany_top_in[73], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[12], chanx_left_in[44], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size9_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_12_sram_inv[0:3]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_0 (
		.bl(bl[0:3]),
		.wl({wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_1 (
		.bl(bl[13:16]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_3 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[5], wl[5], wl[5:6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_5 (
		.bl(bl[1:4]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_7 (
		.bl(bl[5:8]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_9 (
		.bl(bl[9:12]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_11 (
		.bl(bl[13:16]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_13 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[6], wl[6], wl[6:7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_15 (
		.bl(bl[1:4]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_8_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_17 (
		.bl(bl[5:8]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_9_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_19 (
		.bl(bl[9:12]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_10_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_21 (
		.bl(bl[13:16]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_11_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_23 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[7], wl[7], wl[7:8]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_12_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, chany_bottom_in[17], chany_bottom_in[60], chanx_left_in[31], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L1SB_size8_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_0_sram_inv[0:2]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, chany_bottom_in[18], chany_bottom_in[61], chanx_left_in[30], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L1SB_size8_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_1_sram_inv[0:2]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, chany_bottom_in[20], chany_bottom_in[62], chanx_left_in[29], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L1SB_size8_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_2_sram_inv[0:2]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chany_bottom_in[21], chany_bottom_in[64], chanx_left_in[28], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L1SB_size8_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_3_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chany_bottom_in[22], chany_bottom_in[65], chanx_left_in[27], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L1SB_size8_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_4_sram_inv[0:2]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chany_bottom_in[24], chany_bottom_in[66], chanx_left_in[26], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L1SB_size8_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_5_sram_inv[0:2]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chany_bottom_in[25], chany_bottom_in[68], chanx_left_in[25], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L1SB_size8_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_6_sram_inv[0:2]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chany_bottom_in[26], chany_bottom_in[69], chanx_left_in[24], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L1SB_size8_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_7_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chany_bottom_in[28], chany_bottom_in[70], chanx_left_in[23], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L1SB_size8_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_8_sram_inv[0:2]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chany_bottom_in[29], chany_bottom_in[72], chanx_left_in[22], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L1SB_size8_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_9_sram_inv[0:2]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chany_bottom_in[30], chany_bottom_in[73], chanx_left_in[21], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L1SB_size8_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_10_sram_inv[0:2]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_25 (
		.in({chany_top_in[32], chany_top_in[74], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, chanx_left_in[13], chanx_left_in[45], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size8_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_11_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_27 (
		.in({chany_top_in[33], chany_top_in[76], bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, chanx_left_in[14], chanx_left_in[46], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L1SB_size8_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_12_sram_inv[0:2]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_29 (
		.in({chany_top_in[34], chany_top_in[77], bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, chanx_left_in[15], chanx_left_in[47], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L1SB_size8_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_13_sram_inv[0:2]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_2 (
		.bl(bl[4:6]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_4 (
		.bl(bl[7:9]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_1_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_6 (
		.bl(bl[10:12]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_2_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_8 (
		.bl(bl[13:15]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_3_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_10 (
		.bl(bl[16:18]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_4_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_12 (
		.bl({bl[19], bl[0:1]}),
		.wl({wl[0:1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_5_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_14 (
		.bl(bl[2:4]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_6_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_16 (
		.bl(bl[5:7]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_7_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_18 (
		.bl(bl[8:10]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_8_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_20 (
		.bl(bl[11:13]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_9_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_22 (
		.bl(bl[14:16]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_10_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_25 (
		.bl(bl[1:3]),
		.wl({wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_11_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_27 (
		.bl(bl[4:6]),
		.wl({wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_12_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_29 (
		.bl(bl[7:9]),
		.wl({wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_13_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size7 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, chany_bottom_in[32], chany_bottom_in[74], chanx_left_in[20], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L1SB_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size7_0_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_L1SB_size7 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, chany_bottom_in[33], chany_bottom_in[76], chanx_left_in[19], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L1SB_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size7_1_sram_inv[0:2]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_L1SB_size7 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, chany_bottom_in[34], chany_bottom_in[77], chanx_left_in[18], chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L1SB_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size7_2_sram_inv[0:2]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_L1SB_size7 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, chany_bottom_in[36], chany_bottom_in[78], chanx_left_in[17], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L1SB_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size7_3_sram_inv[0:2]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_L1SB_size7 mux_bottom_track_31 (
		.in({chany_top_in[36], chany_top_in[78], bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, chanx_left_in[16], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L1SB_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size7_4_sram_inv[0:2]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_L1SB_size7_mem mem_top_track_24 (
		.bl(bl[17:19]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size7_mem mem_top_track_26 (
		.bl(bl[0:2]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size7_mem mem_top_track_28 (
		.bl(bl[3:5]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size7_mem mem_top_track_30 (
		.bl(bl[6:8]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size7_mem mem_bottom_track_31 (
		.bl(bl[10:12]),
		.wl({wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L1SB_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chany_bottom_in[37], chanx_left_in[16], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_0_sram_inv[0:3]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chany_bottom_in[42], chanx_left_in[12], chanx_left_in[44], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L4SB_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_1_sram_inv[0:3]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chany_bottom_in[44], chanx_left_in[11], chanx_left_in[43], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_2_sram_inv[0:3]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chany_bottom_in[45], chanx_left_in[10], chanx_left_in[42], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L4SB_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_3_sram_inv[0:3]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chany_bottom_in[46], chanx_left_in[9], chanx_left_in[41], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_4_sram_inv[0:3]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chany_bottom_in[53], chanx_left_in[4], chanx_left_in[36], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_5_sram_inv[0:3]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chany_bottom_in[54], chanx_left_in[3], chanx_left_in[35], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_6_sram_inv[0:3]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chany_bottom_in[56], chanx_left_in[2], chanx_left_in[34], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L4SB_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_7_sram_inv[0:3]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_L4SB_size11 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chany_bottom_in[57], chanx_left_in[1], chanx_left_in[33], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_8_sram_inv[0:3]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_33 (
		.in({chany_top_in[37], bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[17], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_9_sram_inv[0:3]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_41 (
		.in({chany_top_in[38], bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[18], chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_10_sram_inv[0:3]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_49 (
		.in({chany_top_in[40], bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[19], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size11_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_11_sram_inv[0:3]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_57 (
		.in({chany_top_in[41], bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[20], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size11_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_12_sram_inv[0:3]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_97 (
		.in({chany_top_in[48], bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_left_in[25], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size11_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_13_sram_inv[0:3]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_105 (
		.in({chany_top_in[49], bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_left_in[26], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L4SB_size11_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_14_sram_inv[0:3]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_113 (
		.in({chany_top_in[50], bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_left_in[27], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size11_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_15_sram_inv[0:3]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_121 (
		.in({chany_top_in[52], bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_left_in[28], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size11_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_16_sram_inv[0:3]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_153 (
		.in({chany_top_in[57], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[0], chanx_left_in[32], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size11_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_17_sram_inv[0:3]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_32 (
		.bl(bl[9:12]),
		.wl({wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_64 (
		.bl(bl[5:8]),
		.wl({wl[3], wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_72 (
		.bl(bl[9:12]),
		.wl({wl[3], wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_80 (
		.bl(bl[13:16]),
		.wl({wl[3], wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_88 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[3], wl[3], wl[3:4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_128 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[4], wl[4], wl[4:5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_136 (
		.bl(bl[1:4]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_144 (
		.bl(bl[5:8]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_top_track_152 (
		.bl(bl[9:12]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_33 (
		.bl(bl[13:16]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_41 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[8], wl[8], wl[8:9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_49 (
		.bl(bl[1:4]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_57 (
		.bl(bl[5:8]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_97 (
		.bl(bl[5:8]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_105 (
		.bl(bl[9:12]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_113 (
		.bl(bl[13:16]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_15_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_121 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[10], wl[10], wl[10:11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_16_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_153 (
		.bl(bl[13:16]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size11_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_17_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chany_bottom_in[38], chanx_left_in[15], chanx_left_in[47], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_0_sram_inv[0:3]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_L4SB_size12 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chany_bottom_in[40], chanx_left_in[14], chanx_left_in[46], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L4SB_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_1_sram_inv[0:3]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_L4SB_size12 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chany_bottom_in[41], chanx_left_in[13], chanx_left_in[45], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L4SB_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_2_sram_inv[0:3]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_L4SB_size12 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_30__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_38__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_46__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_54__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_62__pin_a2f_o_0_, chany_bottom_in[48], chanx_left_in[8], chanx_left_in[40], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_3_sram_inv[0:3]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_L4SB_size12 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_31__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_39__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_47__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_55__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_63__pin_a2f_o_0_, chany_bottom_in[49], chanx_left_in[7], chanx_left_in[39], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_4_sram_inv[0:3]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_L4SB_size12 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_32__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_40__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_48__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_56__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_64__pin_a2f_o_0_, chany_bottom_in[50], chanx_left_in[6], chanx_left_in[38], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L4SB_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_5_sram_inv[0:3]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_L4SB_size12 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_33__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_41__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_49__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_57__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_65__pin_a2f_o_0_, chany_bottom_in[52], chanx_left_in[5], chanx_left_in[37], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_6_sram_inv[0:3]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_L4SB_size12_mem mem_top_track_40 (
		.bl(bl[13:16]),
		.wl({wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_top_track_48 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[2], wl[2], wl[2:3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_top_track_56 (
		.bl(bl[1:4]),
		.wl({wl[3], wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_top_track_96 (
		.bl(bl[1:4]),
		.wl({wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_top_track_104 (
		.bl(bl[5:8]),
		.wl({wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_top_track_112 (
		.bl(bl[9:12]),
		.wl({wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_top_track_120 (
		.bl(bl[13:16]),
		.wl({wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_65 (
		.in({chany_top_in[42], bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[21], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_0_sram_inv[0:3]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_73 (
		.in({chany_top_in[44], bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[22], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_1_sram_inv[0:3]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_81 (
		.in({chany_top_in[45], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[23], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size10_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_2_sram_inv[0:3]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_89 (
		.in({chany_top_in[46], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_left_in[24], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size10_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_3_sram_inv[0:3]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_129 (
		.in({chany_top_in[53], bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_left_in[29], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size10_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_4_sram_inv[0:3]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_137 (
		.in({chany_top_in[54], bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_left_in[30], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L4SB_size10_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_5_sram_inv[0:3]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_145 (
		.in({chany_top_in[56], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_left_in[31], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size10_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_6_sram_inv[0:3]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_65 (
		.bl(bl[9:12]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_73 (
		.bl(bl[13:16]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_81 (
		.bl({bl[17:19], bl[0]}),
		.wl({wl[9], wl[9], wl[9:10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size10_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_89 (
		.bl(bl[1:4]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size10_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_129 (
		.bl(bl[1:4]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size10_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_137 (
		.bl(bl[5:8]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size10_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_145 (
		.bl(bl[9:12]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size10_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_6_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[16], chany_bottom_in[16], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_0_sram_inv[0:1]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_3 (
		.in({chany_top_in[17], chany_bottom_in[0], chany_bottom_in[17], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_1_sram_inv[0:1]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_5 (
		.in({chany_top_in[18], chany_bottom_in[1], chany_bottom_in[18], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_2_sram_inv[0:1]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_7 (
		.in({chany_top_in[20], chany_bottom_in[2], chany_bottom_in[20], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_3_sram_inv[0:1]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_9 (
		.in({chany_top_in[21], chany_bottom_in[3], chany_bottom_in[21], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_4_sram_inv[0:1]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_11 (
		.in({chany_top_in[22], chany_bottom_in[4], chany_bottom_in[22], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_5_sram_inv[0:1]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_13 (
		.in({chany_top_in[24], chany_bottom_in[5], chany_bottom_in[24], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_6_sram_inv[0:1]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_15 (
		.in({chany_top_in[25], chany_bottom_in[6], chany_bottom_in[25], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_7_sram_inv[0:1]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_17 (
		.in({chany_top_in[26], chany_bottom_in[7], chany_bottom_in[26], left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_8_sram_inv[0:1]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_19 (
		.in({chany_top_in[28], chany_bottom_in[8], chany_bottom_in[28], left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_9_sram_inv[0:1]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_21 (
		.in({chany_top_in[29], chany_bottom_in[9], chany_bottom_in[29], left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_10_sram_inv[0:1]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_23 (
		.in({chany_top_in[30], chany_bottom_in[10], chany_bottom_in[30], left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_11_sram_inv[0:1]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_1 (
		.bl(bl[17:18]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_3 (
		.bl({bl[19], bl[0]}),
		.wl(wl[11:12]),
		.mem_out(mux_tree_tapbuf_L1SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_5 (
		.bl(bl[1:2]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_7 (
		.bl(bl[3:4]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_9 (
		.bl(bl[5:6]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_11 (
		.bl(bl[7:8]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_13 (
		.bl(bl[9:10]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_15 (
		.bl(bl[11:12]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_17 (
		.bl(bl[13:14]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_19 (
		.bl(bl[15:16]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_21 (
		.bl(bl[17:18]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_23 (
		.bl({bl[19], bl[0]}),
		.wl(wl[12:13]),
		.mem_out(mux_tree_tapbuf_L1SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3 mux_left_track_25 (
		.in({chany_top_in[32], chany_bottom_in[11], chany_bottom_in[32]}),
		.sram(mux_tree_tapbuf_L1SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_0_sram_inv[0:1]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_L1SB_size3 mux_left_track_27 (
		.in({chany_top_in[33], chany_bottom_in[12], chany_bottom_in[33]}),
		.sram(mux_tree_tapbuf_L1SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_1_sram_inv[0:1]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_L1SB_size3 mux_left_track_29 (
		.in({chany_top_in[34], chany_bottom_in[13], chany_bottom_in[34]}),
		.sram(mux_tree_tapbuf_L1SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_2_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_L1SB_size3 mux_left_track_31 (
		.in({chany_top_in[36], chany_bottom_in[14], chany_bottom_in[36]}),
		.sram(mux_tree_tapbuf_L1SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_3_sram_inv[0:1]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_L1SB_size3_mem mem_left_track_25 (
		.bl(bl[1:2]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_left_track_27 (
		.bl(bl[3:4]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_left_track_29 (
		.bl(bl[5:6]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_left_track_31 (
		.bl(bl[7:8]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_33 (
		.in({chany_top_in[37], chany_bottom_in[15], chany_bottom_in[37], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_35 (
		.in({chany_top_in[38], chany_bottom_in[19], chany_bottom_in[38], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_37 (
		.in({chany_top_in[40], chany_bottom_in[23], chany_bottom_in[40], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_39 (
		.in({chany_top_in[41], chany_bottom_in[27], chany_bottom_in[41], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_49 (
		.in({chany_top_in[48], chany_bottom_in[47:48], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_51 (
		.in({chany_top_in[49], chany_bottom_in[49], chany_bottom_in[51], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_53 (
		.in({chany_top_in[50], chany_bottom_in[50], chany_bottom_in[55], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_55 (
		.in({chany_top_in[52], chany_bottom_in[52], chany_bottom_in[59], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_65 (
		.in({chany_top_in[58], chany_bottom_in[58], chany_bottom_in[79], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_8_sram_inv[0:2]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_33 (
		.bl(bl[9:11]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_35 (
		.bl(bl[12:14]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_37 (
		.bl(bl[15:17]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_39 (
		.bl({bl[18:19], bl[0]}),
		.wl({wl[13], wl[13:14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_49 (
		.bl(bl[9:11]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_51 (
		.bl(bl[12:14]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_53 (
		.bl(bl[15:17]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_55 (
		.bl({bl[18:19], bl[0]}),
		.wl({wl[14], wl[14:15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_65 (
		.bl(bl[9:11]),
		.wl({wl[15], wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_41 (
		.in({chany_top_in[42], chany_bottom_in[31], chany_bottom_in[42], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_0_sram_inv[0:1]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_43 (
		.in({chany_top_in[44], chany_bottom_in[35], chany_bottom_in[44], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_1_sram_inv[0:1]),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_45 (
		.in({chany_top_in[45], chany_bottom_in[39], chany_bottom_in[45], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_2_sram_inv[0:1]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_47 (
		.in({chany_top_in[46], chany_bottom_in[43], chany_bottom_in[46], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_3_sram_inv[0:1]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_57 (
		.in({chany_top_in[53], chany_bottom_in[53], chany_bottom_in[63], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_4_sram_inv[0:1]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_59 (
		.in({chany_top_in[54], chany_bottom_in[54], chany_bottom_in[67], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_5_sram_inv[0:1]),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_61 (
		.in({chany_top_in[56], chany_bottom_in[56], chany_bottom_in[71], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_6_sram_inv[0:1]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_63 (
		.in({chany_top_in[57], chany_bottom_in[57], chany_bottom_in[75], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_7_sram_inv[0:1]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_67 (
		.in({chany_top_in[60], chany_bottom_in[60], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_8_sram_inv[0:1]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_69 (
		.in({chany_top_in[61], chany_bottom_in[61], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_9_sram_inv[0:1]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_71 (
		.in({chany_top_in[62], chany_bottom_in[62], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_10_sram_inv[0:1]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_81 (
		.in({chany_top_in[69], chany_bottom_in[69], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_11_sram_inv[0:1]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_83 (
		.in({chany_top_in[70], chany_bottom_in[70], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_12_sram_inv[0:1]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_85 (
		.in({chany_top_in[72], chany_bottom_in[72], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_13_sram_inv[0:1]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_87 (
		.in({chany_top_in[73], chany_bottom_in[73], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size4_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_14_sram_inv[0:1]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_41 (
		.bl(bl[1:2]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_43 (
		.bl(bl[3:4]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_45 (
		.bl(bl[5:6]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_47 (
		.bl(bl[7:8]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_57 (
		.bl(bl[1:2]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_59 (
		.bl(bl[3:4]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_61 (
		.bl(bl[5:6]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_63 (
		.bl(bl[7:8]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_67 (
		.bl(bl[12:13]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_69 (
		.bl(bl[14:15]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_71 (
		.bl(bl[16:17]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_81 (
		.bl(bl[6:7]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_83 (
		.bl(bl[8:9]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_85 (
		.bl(bl[10:11]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_87 (
		.bl(bl[12:13]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_73 (
		.in({chany_top_in[64], chany_bottom_in[64], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_75 (
		.in({chany_top_in[65], chany_bottom_in[65], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_77 (
		.in({chany_top_in[66], chany_bottom_in[66], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_79 (
		.in({chany_top_in[68], chany_bottom_in[68], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_89 (
		.in({chany_top_in[74], chany_bottom_in[74], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_91 (
		.in({chany_top_in[76], chany_bottom_in[76], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_93 (
		.in({chany_top_in[77], chany_bottom_in[77], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_95 (
		.in({chany_top_in[78], chany_bottom_in[78], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_99 (
		.in({chany_top_in[79], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_101 (
		.in({chany_top_in[75], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_103 (
		.in({chany_top_in[71], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_113 (
		.in({chany_top_in[51], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_115 (
		.in({chany_top_in[47], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_117 (
		.in({chany_top_in[43], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_119 (
		.in({chany_top_in[39], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_129 (
		.in({chany_top_in[19], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_131 (
		.in({chany_top_in[15], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_133 (
		.in({chany_top_in[14], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_135 (
		.in({chany_top_in[13], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_145 (
		.in({chany_top_in[8], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_147 (
		.in({chany_top_in[7], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]),
		.out(chanx_left_out[73]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_149 (
		.in({chany_top_in[6], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]),
		.out(chanx_left_out[74]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_151 (
		.in({chany_top_in[5], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_73 (
		.bl(bl[18:19]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_75 (
		.bl(bl[0:1]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_77 (
		.bl(bl[2:3]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_79 (
		.bl(bl[4:5]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_89 (
		.bl(bl[14:15]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_91 (
		.bl(bl[16:17]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_93 (
		.bl(bl[18:19]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_95 (
		.bl(bl[0:1]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_99 (
		.bl(bl[3:4]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_101 (
		.bl(bl[5:6]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_103 (
		.bl(bl[7:8]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_113 (
		.bl(bl[13:14]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_115 (
		.bl(bl[15:16]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_117 (
		.bl(bl[17:18]),
		.wl({wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_119 (
		.bl({bl[19], bl[0]}),
		.wl(wl[17:18]),
		.mem_out(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_129 (
		.bl(bl[5:6]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_131 (
		.bl(bl[7:8]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_133 (
		.bl(bl[9:10]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_135 (
		.bl(bl[11:12]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_145 (
		.bl(bl[17:18]),
		.wl({wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_147 (
		.bl({bl[19], bl[0]}),
		.wl(wl[18:19]),
		.mem_out(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_149 (
		.bl(bl[1:2]),
		.wl({wl[19], wl[19]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_151 (
		.bl(bl[3:4]),
		.wl({wl[19], wl[19]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_97 (
		.in({left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_0_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_0_sram_inv),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_105 (
		.in({chany_top_in[67], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_1_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_1_sram_inv),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_107 (
		.in({chany_top_in[63], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_2_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_2_sram_inv),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_109 (
		.in({chany_top_in[59], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_3_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_3_sram_inv),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_111 (
		.in({chany_top_in[55], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_4_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_4_sram_inv),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_121 (
		.in({chany_top_in[35], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_5_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_5_sram_inv),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_123 (
		.in({chany_top_in[31], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_6_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_6_sram_inv),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_125 (
		.in({chany_top_in[27], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_7_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_7_sram_inv),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_127 (
		.in({chany_top_in[23], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_8_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_8_sram_inv),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_137 (
		.in({chany_top_in[12], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_9_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_9_sram_inv),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_139 (
		.in({chany_top_in[11], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_10_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_10_sram_inv),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_141 (
		.in({chany_top_in[10], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_11_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_11_sram_inv),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_143 (
		.in({chany_top_in[9], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_12_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_12_sram_inv),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_153 (
		.in({chany_top_in[4], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_13_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_13_sram_inv),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_155 (
		.in({chany_top_in[3], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_14_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_14_sram_inv),
		.out(chanx_left_out[77]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_157 (
		.in({chany_top_in[2], left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_15_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_15_sram_inv),
		.out(chanx_left_out[78]));

	mux_tree_tapbuf_L4SB_size2 mux_left_track_159 (
		.in({chany_top_in[1], left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_16_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_16_sram_inv),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_97 (
		.bl(bl[2]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_0_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_0_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_105 (
		.bl(bl[9]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_1_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_1_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_107 (
		.bl(bl[10]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_2_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_2_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_109 (
		.bl(bl[11]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_3_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_3_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_111 (
		.bl(bl[12]),
		.wl(wl[17]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_4_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_4_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_121 (
		.bl(bl[1]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_5_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_5_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_123 (
		.bl(bl[2]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_6_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_6_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_125 (
		.bl(bl[3]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_7_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_7_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_127 (
		.bl(bl[4]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_8_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_8_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_137 (
		.bl(bl[13]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_9_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_9_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_139 (
		.bl(bl[14]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_10_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_10_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_141 (
		.bl(bl[15]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_11_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_11_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_143 (
		.bl(bl[16]),
		.wl(wl[18]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_12_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_12_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_153 (
		.bl(bl[5]),
		.wl(wl[19]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_13_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_13_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_155 (
		.bl(bl[6]),
		.wl(wl[19]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_14_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_14_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_157 (
		.bl(bl[7]),
		.wl(wl[19]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_15_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_15_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_left_track_159 (
		.bl(bl[8]),
		.wl(wl[19]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_16_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_16_sram_inv));

endmodule
// ----- END Verilog module for sb_10__1_ -----

//----- Default net type -----
`default_nettype none



