//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_1__0_ -----
module sb_1__0_(chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                chanx_right_in,
                chanx_left_in,
                bl,
                wl,
                chany_top_out,
                chanx_right_out,
                chanx_left_out);
//----- INPUT PORTS -----
input [0:79] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:79] chanx_right_in;
//----- INPUT PORTS -----
input [0:79] chanx_left_in;
//----- INPUT PORTS -----
input [0:17] bl;
//----- INPUT PORTS -----
input [0:16] wl;
//----- OUTPUT PORTS -----
output [0:79] chany_top_out;
//----- OUTPUT PORTS -----
output [0:79] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:79] chanx_left_out;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_L1SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_12_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_13_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_14_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_15_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_16_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_17_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_18_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_19_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_20_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_21_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_22_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_23_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_24_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_25_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_26_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_10_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_11_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_12_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_13_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_14_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_15_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_16_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_6_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_7_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_8_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_9_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_30_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_31_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_32_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_33_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_34_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_35_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_36_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_37_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_38_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_39_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_40_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_17_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_18_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_19_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_20_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_21_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_22_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_23_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_24_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_25_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_26_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_27_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_27_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_28_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_28_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_29_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_29_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_30_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_30_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L1SB_size5 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, chanx_right_in[1], chanx_right_in[16], chanx_left_in[0], chanx_left_in[16]}),
		.sram(mux_tree_tapbuf_L1SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[32], chany_top_in[64], chanx_left_in[17], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L1SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_1_sram_inv[0:2]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[33], chany_top_in[65], chanx_left_in[18], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L1SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_2_sram_inv[0:2]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[34], chany_top_in[66], chanx_left_in[20], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L1SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_3_sram_inv[0:2]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_8 (
		.in({chany_top_in[3], chany_top_in[35], chany_top_in[67], chanx_left_in[21], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L1SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_4_sram_inv[0:2]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_10 (
		.in({chany_top_in[4], chany_top_in[36], chany_top_in[68], chanx_left_in[22], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L1SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_5_sram_inv[0:2]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_12 (
		.in({chany_top_in[5], chany_top_in[37], chany_top_in[69], chanx_left_in[24], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L1SB_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_6_sram_inv[0:2]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_14 (
		.in({chany_top_in[6], chany_top_in[38], chany_top_in[70], chanx_left_in[25], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L1SB_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_7_sram_inv[0:2]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_16 (
		.in({chany_top_in[7], chany_top_in[39], chany_top_in[71], chanx_left_in[26], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L1SB_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_8_sram_inv[0:2]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_18 (
		.in({chany_top_in[8], chany_top_in[40], chany_top_in[72], chanx_left_in[28], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L1SB_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_9_sram_inv[0:2]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_20 (
		.in({chany_top_in[9], chany_top_in[41], chany_top_in[73], chanx_left_in[29], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_10_sram_inv[0:2]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_22 (
		.in({chany_top_in[10], chany_top_in[42], chany_top_in[74], chanx_left_in[30], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_11_sram_inv[0:2]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_24 (
		.in({chany_top_in[11], chany_top_in[43], chany_top_in[75], chanx_left_in[32], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L1SB_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_12_sram_inv[0:2]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_26 (
		.in({chany_top_in[12], chany_top_in[44], chany_top_in[76], chanx_left_in[33], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_13_sram_inv[0:2]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_28 (
		.in({chany_top_in[13], chany_top_in[45], chany_top_in[77], chanx_left_in[34], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_14_sram_inv[0:2]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_30 (
		.in({chany_top_in[14], chany_top_in[46], chany_top_in[78], chanx_left_in[36], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L1SB_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_15_sram_inv[0:2]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_L1SB_size5 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[32], chany_top_in[64], chanx_right_in[16], chanx_right_in[58]}),
		.sram(mux_tree_tapbuf_L1SB_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_16_sram_inv[0:2]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_L1SB_size5_mem mem_top_track_0 (
		.bl(bl[0:2]),
		.wl({wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_2 (
		.bl(bl[11:13]),
		.wl({wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_4 (
		.bl(bl[14:16]),
		.wl({wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_6 (
		.bl({bl[17], bl[0:1]}),
		.wl({wl[8:9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_8 (
		.bl(bl[2:4]),
		.wl({wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_10 (
		.bl(bl[5:7]),
		.wl({wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_12 (
		.bl(bl[8:10]),
		.wl({wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_14 (
		.bl(bl[11:13]),
		.wl({wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_16 (
		.bl(bl[14:16]),
		.wl({wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_18 (
		.bl({bl[17], bl[0:1]}),
		.wl({wl[9:10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_20 (
		.bl(bl[2:4]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_22 (
		.bl(bl[5:7]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_24 (
		.bl(bl[8:10]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_26 (
		.bl(bl[11:13]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_28 (
		.bl(bl[14:16]),
		.wl({wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_30 (
		.bl({bl[17], bl[0:1]}),
		.wl({wl[10:11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_left_track_1 (
		.bl({bl[16:17], bl[0]}),
		.wl({wl[12], wl[12:13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, chanx_right_in[2], chanx_right_in[17], chanx_left_in[17]}),
		.sram(mux_tree_tapbuf_L1SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_0_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, chanx_right_in[3], chanx_right_in[18], chanx_left_in[18]}),
		.sram(mux_tree_tapbuf_L1SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_1_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, chanx_right_in[4], chanx_right_in[20], chanx_left_in[20]}),
		.sram(mux_tree_tapbuf_L1SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_2_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_right_in[5], chanx_right_in[21], chanx_left_in[21]}),
		.sram(mux_tree_tapbuf_L1SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_3_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_right_in[6], chanx_right_in[22], chanx_left_in[22]}),
		.sram(mux_tree_tapbuf_L1SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_4_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_right_in[7], chanx_right_in[24], chanx_left_in[24]}),
		.sram(mux_tree_tapbuf_L1SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_5_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[8], chanx_right_in[25], chanx_left_in[25]}),
		.sram(mux_tree_tapbuf_L1SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_6_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_right_in[9], chanx_right_in[26], chanx_left_in[26]}),
		.sram(mux_tree_tapbuf_L1SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_7_sram_inv[0:1]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_right_in[10], chanx_right_in[28], chanx_left_in[28]}),
		.sram(mux_tree_tapbuf_L1SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_8_sram_inv[0:1]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_right_in[11], chanx_right_in[29], chanx_left_in[29]}),
		.sram(mux_tree_tapbuf_L1SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_9_sram_inv[0:1]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_L1SB_size4 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_right_in[12], chanx_right_in[30], chanx_left_in[30]}),
		.sram(mux_tree_tapbuf_L1SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_10_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_L1SB_size4 mux_right_track_0 (
		.in({chany_top_in[31], chany_top_in[63], chanx_left_in[16], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L1SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_11_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_3 (
		.in({chany_top_in[31], chany_top_in[63], chanx_right_in[17], chanx_right_in[60]}),
		.sram(mux_tree_tapbuf_L1SB_size4_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_12_sram_inv[0:1]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_5 (
		.in({chany_top_in[30], chany_top_in[62], chanx_right_in[18], chanx_right_in[61]}),
		.sram(mux_tree_tapbuf_L1SB_size4_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_13_sram_inv[0:1]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_7 (
		.in({chany_top_in[29], chany_top_in[61], chanx_right_in[20], chanx_right_in[62]}),
		.sram(mux_tree_tapbuf_L1SB_size4_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_14_sram_inv[0:1]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_9 (
		.in({chany_top_in[28], chany_top_in[60], chanx_right_in[21], chanx_right_in[64]}),
		.sram(mux_tree_tapbuf_L1SB_size4_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_15_sram_inv[0:1]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_11 (
		.in({chany_top_in[27], chany_top_in[59], chanx_right_in[22], chanx_right_in[65]}),
		.sram(mux_tree_tapbuf_L1SB_size4_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_16_sram_inv[0:1]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_13 (
		.in({chany_top_in[26], chany_top_in[58], chanx_right_in[24], chanx_right_in[66]}),
		.sram(mux_tree_tapbuf_L1SB_size4_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_17_sram_inv[0:1]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_15 (
		.in({chany_top_in[25], chany_top_in[57], chanx_right_in[25], chanx_right_in[68]}),
		.sram(mux_tree_tapbuf_L1SB_size4_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_18_sram_inv[0:1]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_17 (
		.in({chany_top_in[24], chany_top_in[56], chanx_right_in[26], chanx_right_in[69]}),
		.sram(mux_tree_tapbuf_L1SB_size4_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_19_sram_inv[0:1]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_19 (
		.in({chany_top_in[23], chany_top_in[55], chanx_right_in[28], chanx_right_in[70]}),
		.sram(mux_tree_tapbuf_L1SB_size4_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_20_sram_inv[0:1]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_21 (
		.in({chany_top_in[22], chany_top_in[54], chanx_right_in[29], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size4_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_21_sram_inv[0:1]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_23 (
		.in({chany_top_in[21], chany_top_in[53], chanx_right_in[30], chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size4_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_22_sram_inv[0:1]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_25 (
		.in({chany_top_in[20], chany_top_in[52], chanx_right_in[32], chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_L1SB_size4_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_23_sram_inv[0:1]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_27 (
		.in({chany_top_in[19], chany_top_in[51], chanx_right_in[33], chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size4_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_24_sram_inv[0:1]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_29 (
		.in({chany_top_in[18], chany_top_in[50], chanx_right_in[34], chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size4_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_25_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_31 (
		.in({chany_top_in[17], chany_top_in[49], chanx_right_in[36], chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_L1SB_size4_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_26_sram_inv[0:1]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_2 (
		.bl(bl[3:4]),
		.wl({wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_4 (
		.bl(bl[5:6]),
		.wl({wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_6 (
		.bl(bl[7:8]),
		.wl({wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_8 (
		.bl(bl[9:10]),
		.wl({wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_10 (
		.bl(bl[11:12]),
		.wl({wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_12 (
		.bl(bl[13:14]),
		.wl({wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_14 (
		.bl(bl[15:16]),
		.wl({wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_16 (
		.bl({bl[17], bl[0]}),
		.wl(wl[0:1]),
		.mem_out(mux_tree_tapbuf_L1SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_18 (
		.bl(bl[1:2]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_20 (
		.bl(bl[3:4]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_22 (
		.bl(bl[5:6]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_right_track_0 (
		.bl(bl[9:10]),
		.wl({wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_3 (
		.bl(bl[1:2]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_12_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_5 (
		.bl(bl[3:4]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_13_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_7 (
		.bl(bl[5:6]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_14_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_9 (
		.bl(bl[7:8]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_15_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_11 (
		.bl(bl[9:10]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_16_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_13 (
		.bl(bl[11:12]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_17_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_15 (
		.bl(bl[13:14]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_18_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_17 (
		.bl(bl[15:16]),
		.wl({wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_19_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_19 (
		.bl({bl[17], bl[0]}),
		.wl(wl[13:14]),
		.mem_out(mux_tree_tapbuf_L1SB_size4_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_20_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_21 (
		.bl(bl[1:2]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_21_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_23 (
		.bl(bl[3:4]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_22_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_25 (
		.bl(bl[5:6]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_23_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_27 (
		.bl(bl[7:8]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_24_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_29 (
		.bl(bl[9:10]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_25_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_31 (
		.bl(bl[11:12]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L1SB_size4_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_26_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_24 (
		.in({chanx_right_in[13], chanx_right_in[32], chanx_left_in[32]}),
		.sram(mux_tree_tapbuf_L1SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_0_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_26 (
		.in({chanx_right_in[14], chanx_right_in[33], chanx_left_in[33]}),
		.sram(mux_tree_tapbuf_L1SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_1_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_28 (
		.in({chanx_right_in[15], chanx_right_in[34], chanx_left_in[34]}),
		.sram(mux_tree_tapbuf_L1SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_2_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_30 (
		.in({chanx_right_in[19], chanx_right_in[36], chanx_left_in[36]}),
		.sram(mux_tree_tapbuf_L1SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_3_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_24 (
		.bl(bl[7:8]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_26 (
		.bl(bl[9:10]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_28 (
		.bl(bl[11:12]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_30 (
		.bl(bl[13:14]),
		.wl({wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_right_in[23], chanx_right_in[37], chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_34 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_right_in[27], chanx_right_in[38], chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]),
		.out(chany_top_out[17]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_right_in[31], chanx_right_in[40], chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]),
		.out(chany_top_out[18]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_right_in[35], chanx_right_in[41], chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]),
		.out(chany_top_out[19]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_right_in[48], chanx_right_in[55], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_right_in[49], chanx_right_in[59], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]),
		.out(chany_top_out[25]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_52 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_right_in[50], chanx_right_in[63], chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]),
		.out(chany_top_out[26]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_54 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_right_in[52], chanx_right_in[67], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]),
		.out(chany_top_out[27]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_32 (
		.bl(bl[15:17]),
		.wl({wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_34 (
		.bl(bl[0:2]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_36 (
		.bl(bl[3:5]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_38 (
		.bl(bl[6:8]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_48 (
		.bl({bl[17], bl[0:1]}),
		.wl({wl[2:3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_50 (
		.bl(bl[2:4]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_52 (
		.bl(bl[5:7]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_54 (
		.bl(bl[8:10]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_right_in[39], chanx_right_in[42], chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_0_sram_inv[0:1]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_right_in[43:44], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_1_sram_inv[0:1]),
		.out(chany_top_out[21]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_right_in[45], chanx_right_in[47], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_2_sram_inv[0:1]),
		.out(chany_top_out[22]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_46 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[46], chanx_right_in[51], chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_3_sram_inv[0:1]),
		.out(chany_top_out[23]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_right_in[53], chanx_right_in[71], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_4_sram_inv[0:1]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_right_in[54], chanx_right_in[75], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_5_sram_inv[0:1]),
		.out(chany_top_out[29]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_right_in[56], chanx_right_in[79], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_6_sram_inv[0:1]),
		.out(chany_top_out[30]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_right_in[58], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L4SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_7_sram_inv[0:1]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_right_in[60], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_8_sram_inv[0:1]),
		.out(chany_top_out[33]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_right_in[61], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_9_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_70 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_right_in[62], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L4SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_10_sram_inv[0:1]),
		.out(chany_top_out[35]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_right_in[69], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_11_sram_inv[0:1]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_right_in[70], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L4SB_size4_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_12_sram_inv[0:1]),
		.out(chany_top_out[41]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_right_in[72], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size4_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_13_sram_inv[0:1]),
		.out(chany_top_out[42]));

	mux_tree_tapbuf_L4SB_size4 mux_top_track_86 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_right_in[73], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size4_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_14_sram_inv[0:1]),
		.out(chany_top_out[43]));

	mux_tree_tapbuf_L4SB_size4 mux_right_track_32 (
		.in({chany_top_in[15], chany_top_in[47], chany_top_in[79], chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size4_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_15_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_41 (
		.in({chany_top_in[15], chany_top_in[47], chany_top_in[79], chanx_right_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size4_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_16_sram_inv[0:1]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_49 (
		.in({chany_top_in[14], chany_top_in[46], chany_top_in[78], chanx_right_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size4_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_17_sram_inv[0:1]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_57 (
		.in({chany_top_in[13], chany_top_in[45], chany_top_in[77], chanx_right_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size4_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_18_sram_inv[0:1]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_65 (
		.in({chany_top_in[12], chany_top_in[44], chany_top_in[76], chanx_right_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size4_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_19_sram_inv[0:1]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_73 (
		.in({chany_top_in[11], chany_top_in[43], chany_top_in[75], chanx_right_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size4_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_20_sram_inv[0:1]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_81 (
		.in({chany_top_in[10], chany_top_in[42], chany_top_in[74], chanx_right_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size4_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_21_sram_inv[0:1]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_89 (
		.in({chany_top_in[9], chany_top_in[41], chany_top_in[73], chanx_right_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size4_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_22_sram_inv[0:1]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_97 (
		.in({chany_top_in[8], chany_top_in[40], chany_top_in[72], chanx_right_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size4_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_23_sram_inv[0:1]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_105 (
		.in({chany_top_in[7], chany_top_in[39], chany_top_in[71], chanx_right_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size4_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_24_sram_inv[0:1]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_113 (
		.in({chany_top_in[6], chany_top_in[38], chany_top_in[70], chanx_right_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size4_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_25_sram_inv[0:1]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_121 (
		.in({chany_top_in[5], chany_top_in[37], chany_top_in[69], chanx_right_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size4_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_26_sram_inv[0:1]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_129 (
		.in({chany_top_in[4], chany_top_in[36], chany_top_in[68], chanx_right_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size4_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_27_sram_inv[0:1]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_137 (
		.in({chany_top_in[3], chany_top_in[35], chany_top_in[67], chanx_right_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size4_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_28_sram_inv[0:1]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_145 (
		.in({chany_top_in[2], chany_top_in[34], chany_top_in[66], chanx_right_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size4_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_29_sram_inv[0:1]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_153 (
		.in({chany_top_in[1], chany_top_in[33], chany_top_in[65], chanx_right_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size4_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_30_sram_inv[0:1]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_40 (
		.bl(bl[9:10]),
		.wl({wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_42 (
		.bl(bl[11:12]),
		.wl({wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_44 (
		.bl(bl[13:14]),
		.wl({wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_46 (
		.bl(bl[15:16]),
		.wl({wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_56 (
		.bl(bl[11:12]),
		.wl({wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_58 (
		.bl(bl[13:14]),
		.wl({wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_60 (
		.bl(bl[15:16]),
		.wl({wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_64 (
		.bl(bl[1:2]),
		.wl({wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_66 (
		.bl(bl[3:4]),
		.wl({wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_68 (
		.bl(bl[5:6]),
		.wl({wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_70 (
		.bl(bl[7:8]),
		.wl({wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_80 (
		.bl({bl[17], bl[0]}),
		.wl(wl[4:5]),
		.mem_out(mux_tree_tapbuf_L4SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_82 (
		.bl(bl[1:2]),
		.wl({wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_84 (
		.bl(bl[3:4]),
		.wl({wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_top_track_86 (
		.bl(bl[5:6]),
		.wl({wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_right_track_32 (
		.bl(bl[2:3]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_41 (
		.bl(bl[15:16]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_16_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_49 (
		.bl({bl[17], bl[0]}),
		.wl(wl[14:15]),
		.mem_out(mux_tree_tapbuf_L4SB_size4_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_17_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_57 (
		.bl(bl[1:2]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_65 (
		.bl(bl[3:4]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_19_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_73 (
		.bl(bl[5:6]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_20_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_81 (
		.bl(bl[7:8]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_21_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_89 (
		.bl(bl[9:10]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_22_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_97 (
		.bl(bl[11:12]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_23_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_105 (
		.bl(bl[13:14]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_24_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_113 (
		.bl(bl[15:16]),
		.wl({wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_25_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_121 (
		.bl({bl[17], bl[0]}),
		.wl(wl[15:16]),
		.mem_out(mux_tree_tapbuf_L4SB_size4_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_26_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_129 (
		.bl(bl[1:2]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_27_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_137 (
		.bl(bl[3:4]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_28_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_145 (
		.bl(bl[5:6]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_29_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_153 (
		.bl(bl[7:8]),
		.wl({wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L4SB_size4_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_30_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_62 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[57], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]),
		.out(chany_top_out[31]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_right_in[64], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_right_in[65], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]),
		.out(chany_top_out[37]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_right_in[66], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]),
		.out(chany_top_out[38]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_78 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[68], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]),
		.out(chany_top_out[39]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_right_in[74], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_right_in[76], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]),
		.out(chany_top_out[45]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_right_in[77], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]),
		.out(chany_top_out[46]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_94 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[78], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]),
		.out(chany_top_out[47]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]),
		.out(chany_top_out[49]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]),
		.out(chany_top_out[50]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_102 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]),
		.out(chany_top_out[51]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]),
		.out(chany_top_out[57]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]),
		.out(chany_top_out[58]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_118 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[39]}),
		.sram(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]),
		.out(chany_top_out[59]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[19]}),
		.sram(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[15]}),
		.sram(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]),
		.out(chany_top_out[65]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[14]}),
		.sram(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]),
		.out(chany_top_out[66]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_134 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[13]}),
		.sram(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]),
		.out(chany_top_out[67]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[8]}),
		.sram(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[7]}),
		.sram(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]),
		.out(chany_top_out[73]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[6]}),
		.sram(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]),
		.out(chany_top_out[74]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_150 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[5]}),
		.sram(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]),
		.out(chany_top_out[75]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_158 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[0], chanx_left_in[1]}),
		.sram(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]),
		.out(chany_top_out[79]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_40 (
		.in({chany_top_in[16], chany_top_in[48], chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_48 (
		.in({chany_top_in[17], chany_top_in[49], chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_56 (
		.in({chany_top_in[18], chany_top_in[50], chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_64 (
		.in({chany_top_in[19], chany_top_in[51], chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_72 (
		.in({chany_top_in[20], chany_top_in[52], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_80 (
		.in({chany_top_in[21], chany_top_in[53], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_30_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_88 (
		.in({chany_top_in[22], chany_top_in[54], chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_31_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_96 (
		.in({chany_top_in[23], chany_top_in[55], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_32_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_104 (
		.in({chany_top_in[24], chany_top_in[56], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_33_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_112 (
		.in({chany_top_in[25], chany_top_in[57], chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_34_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_120 (
		.in({chany_top_in[26], chany_top_in[58], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_35_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_128 (
		.in({chany_top_in[27], chany_top_in[59], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_36_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_136 (
		.in({chany_top_in[28], chany_top_in[60], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_37_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_144 (
		.in({chany_top_in[29], chany_top_in[61], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_38_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_152 (
		.in({chany_top_in[30], chany_top_in[62], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_39_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_33 (
		.in({chany_top_in[16], chany_top_in[48], chanx_right_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_40_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_62 (
		.bl({bl[17], bl[0]}),
		.wl(wl[3:4]),
		.mem_out(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_72 (
		.bl(bl[9:10]),
		.wl({wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_74 (
		.bl(bl[11:12]),
		.wl({wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_76 (
		.bl(bl[13:14]),
		.wl({wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_78 (
		.bl(bl[15:16]),
		.wl({wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_88 (
		.bl(bl[7:8]),
		.wl({wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_90 (
		.bl(bl[9:10]),
		.wl({wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_92 (
		.bl(bl[11:12]),
		.wl({wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_94 (
		.bl(bl[13:14]),
		.wl({wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_98 (
		.bl(bl[16:17]),
		.wl({wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_100 (
		.bl(bl[0:1]),
		.wl({wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_102 (
		.bl(bl[2:3]),
		.wl({wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_112 (
		.bl(bl[8:9]),
		.wl({wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_114 (
		.bl(bl[10:11]),
		.wl({wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_116 (
		.bl(bl[12:13]),
		.wl({wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_118 (
		.bl(bl[14:15]),
		.wl({wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_128 (
		.bl(bl[2:3]),
		.wl({wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_130 (
		.bl(bl[4:5]),
		.wl({wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_132 (
		.bl(bl[6:7]),
		.wl({wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_134 (
		.bl(bl[8:9]),
		.wl({wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_144 (
		.bl(bl[14:15]),
		.wl({wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_146 (
		.bl(bl[16:17]),
		.wl({wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_148 (
		.bl(bl[0:1]),
		.wl({wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_150 (
		.bl(bl[2:3]),
		.wl({wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_158 (
		.bl(bl[7:8]),
		.wl({wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_40 (
		.bl(bl[4:5]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_48 (
		.bl(bl[6:7]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_56 (
		.bl(bl[8:9]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_64 (
		.bl(bl[10:11]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_72 (
		.bl(bl[12:13]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_80 (
		.bl(bl[14:15]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_88 (
		.bl(bl[16:17]),
		.wl({wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_96 (
		.bl(bl[0:1]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_104 (
		.bl(bl[2:3]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_112 (
		.bl(bl[4:5]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_120 (
		.bl(bl[6:7]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_128 (
		.bl(bl[8:9]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_136 (
		.bl(bl[10:11]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_144 (
		.bl(bl[12:13]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_152 (
		.bl(bl[14:15]),
		.wl({wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_33 (
		.bl(bl[13:14]),
		.wl({wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_0_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_0_sram_inv),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size2_1_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_1_sram_inv),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_106 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size2_2_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_2_sram_inv),
		.out(chany_top_out[53]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size2_3_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_3_sram_inv),
		.out(chany_top_out[54]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_110 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size2_4_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_4_sram_inv),
		.out(chany_top_out[55]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_left_in[35]}),
		.sram(mux_tree_tapbuf_L4SB_size2_5_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_5_sram_inv),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[31]}),
		.sram(mux_tree_tapbuf_L4SB_size2_6_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_6_sram_inv),
		.out(chany_top_out[61]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_124 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[27]}),
		.sram(mux_tree_tapbuf_L4SB_size2_7_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_7_sram_inv),
		.out(chany_top_out[62]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_126 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[23]}),
		.sram(mux_tree_tapbuf_L4SB_size2_8_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_8_sram_inv),
		.out(chany_top_out[63]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_left_in[12]}),
		.sram(mux_tree_tapbuf_L4SB_size2_9_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_9_sram_inv),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[11]}),
		.sram(mux_tree_tapbuf_L4SB_size2_10_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_10_sram_inv),
		.out(chany_top_out[69]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[10]}),
		.sram(mux_tree_tapbuf_L4SB_size2_11_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_11_sram_inv),
		.out(chany_top_out[70]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_142 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[9]}),
		.sram(mux_tree_tapbuf_L4SB_size2_12_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_12_sram_inv),
		.out(chany_top_out[71]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_left_in[4]}),
		.sram(mux_tree_tapbuf_L4SB_size2_13_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_13_sram_inv),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[3]}),
		.sram(mux_tree_tapbuf_L4SB_size2_14_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_14_sram_inv),
		.out(chany_top_out[77]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[2]}),
		.sram(mux_tree_tapbuf_L4SB_size2_15_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_15_sram_inv),
		.out(chany_top_out[78]));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_96 (
		.bl(bl[15]),
		.wl(wl[5]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_0_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_0_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_104 (
		.bl(bl[4]),
		.wl(wl[6]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_1_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_1_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_106 (
		.bl(bl[5]),
		.wl(wl[6]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_2_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_2_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_108 (
		.bl(bl[6]),
		.wl(wl[6]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_3_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_3_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_110 (
		.bl(bl[7]),
		.wl(wl[6]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_4_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_4_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_120 (
		.bl(bl[16]),
		.wl(wl[6]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_5_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_5_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_122 (
		.bl(bl[17]),
		.wl(wl[6]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_6_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_6_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_124 (
		.bl(bl[0]),
		.wl(wl[7]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_7_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_7_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_126 (
		.bl(bl[1]),
		.wl(wl[7]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_8_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_8_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_136 (
		.bl(bl[10]),
		.wl(wl[7]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_9_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_9_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_138 (
		.bl(bl[11]),
		.wl(wl[7]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_10_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_10_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_140 (
		.bl(bl[12]),
		.wl(wl[7]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_11_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_11_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_142 (
		.bl(bl[13]),
		.wl(wl[7]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_12_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_12_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_152 (
		.bl(bl[4]),
		.wl(wl[8]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_13_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_13_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_154 (
		.bl(bl[5]),
		.wl(wl[8]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_14_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_14_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_156 (
		.bl(bl[6]),
		.wl(wl[8]),
		.mem_out(mux_tree_tapbuf_L4SB_size2_15_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_15_sram_inv));

endmodule
// ----- END Verilog module for sb_1__0_ -----

//----- Default net type -----
`default_nettype none



