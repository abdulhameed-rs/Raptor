//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Connection Blocks[1][1]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for cbx_1__1_ -----
module cbx_1__1_(chanx_left_in,
                 chanx_right_in,
                 bl,
                 wl,
                 chanx_left_out,
                 chanx_right_out,
                 bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_20__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_21__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_22__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_23__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_24__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_25__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_26__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_27__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_28__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_29__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_30__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_31__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_32__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_33__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_34__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_35__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_36__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_37__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_38__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_39__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_40__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_41__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_42__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_43__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_44__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_45__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_46__pin_f2a_i_0_,
                 bottom_grid_top_width_0_height_0_subtile_47__pin_f2a_i_0_);
//----- INPUT PORTS -----
input [0:79] chanx_left_in;
//----- INPUT PORTS -----
input [0:79] chanx_right_in;
//----- INPUT PORTS -----
input [0:15] bl;
//----- INPUT PORTS -----
input [0:14] wl;
//----- OUTPUT PORTS -----
output [0:79] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:79] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_20__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_21__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_22__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_23__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_24__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_25__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_26__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_27__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_28__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_29__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_30__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_31__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_32__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_33__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_34__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_35__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_36__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_37__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_38__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_39__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_40__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_41__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_42__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_43__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_44__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_45__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_46__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_grid_top_width_0_height_0_subtile_47__pin_f2a_i_0_;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:4] mux_tree_tapbuf_size18_0_sram;
wire [0:4] mux_tree_tapbuf_size18_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_10_sram;
wire [0:4] mux_tree_tapbuf_size18_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_11_sram;
wire [0:4] mux_tree_tapbuf_size18_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_12_sram;
wire [0:4] mux_tree_tapbuf_size18_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_13_sram;
wire [0:4] mux_tree_tapbuf_size18_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_14_sram;
wire [0:4] mux_tree_tapbuf_size18_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_15_sram;
wire [0:4] mux_tree_tapbuf_size18_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_16_sram;
wire [0:4] mux_tree_tapbuf_size18_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_17_sram;
wire [0:4] mux_tree_tapbuf_size18_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_18_sram;
wire [0:4] mux_tree_tapbuf_size18_18_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_19_sram;
wire [0:4] mux_tree_tapbuf_size18_19_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_1_sram;
wire [0:4] mux_tree_tapbuf_size18_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_20_sram;
wire [0:4] mux_tree_tapbuf_size18_20_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_21_sram;
wire [0:4] mux_tree_tapbuf_size18_21_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_22_sram;
wire [0:4] mux_tree_tapbuf_size18_22_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_23_sram;
wire [0:4] mux_tree_tapbuf_size18_23_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_24_sram;
wire [0:4] mux_tree_tapbuf_size18_24_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_25_sram;
wire [0:4] mux_tree_tapbuf_size18_25_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_26_sram;
wire [0:4] mux_tree_tapbuf_size18_26_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_27_sram;
wire [0:4] mux_tree_tapbuf_size18_27_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_28_sram;
wire [0:4] mux_tree_tapbuf_size18_28_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_29_sram;
wire [0:4] mux_tree_tapbuf_size18_29_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_2_sram;
wire [0:4] mux_tree_tapbuf_size18_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_30_sram;
wire [0:4] mux_tree_tapbuf_size18_30_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_31_sram;
wire [0:4] mux_tree_tapbuf_size18_31_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_32_sram;
wire [0:4] mux_tree_tapbuf_size18_32_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_33_sram;
wire [0:4] mux_tree_tapbuf_size18_33_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_34_sram;
wire [0:4] mux_tree_tapbuf_size18_34_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_35_sram;
wire [0:4] mux_tree_tapbuf_size18_35_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_36_sram;
wire [0:4] mux_tree_tapbuf_size18_36_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_37_sram;
wire [0:4] mux_tree_tapbuf_size18_37_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_38_sram;
wire [0:4] mux_tree_tapbuf_size18_38_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_39_sram;
wire [0:4] mux_tree_tapbuf_size18_39_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_3_sram;
wire [0:4] mux_tree_tapbuf_size18_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_40_sram;
wire [0:4] mux_tree_tapbuf_size18_40_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_41_sram;
wire [0:4] mux_tree_tapbuf_size18_41_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_42_sram;
wire [0:4] mux_tree_tapbuf_size18_42_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_43_sram;
wire [0:4] mux_tree_tapbuf_size18_43_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_44_sram;
wire [0:4] mux_tree_tapbuf_size18_44_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_45_sram;
wire [0:4] mux_tree_tapbuf_size18_45_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_46_sram;
wire [0:4] mux_tree_tapbuf_size18_46_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_47_sram;
wire [0:4] mux_tree_tapbuf_size18_47_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_4_sram;
wire [0:4] mux_tree_tapbuf_size18_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_5_sram;
wire [0:4] mux_tree_tapbuf_size18_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_6_sram;
wire [0:4] mux_tree_tapbuf_size18_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_7_sram;
wire [0:4] mux_tree_tapbuf_size18_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_8_sram;
wire [0:4] mux_tree_tapbuf_size18_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_9_sram;
wire [0:4] mux_tree_tapbuf_size18_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[0] = chanx_left_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[1] = chanx_left_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[2] = chanx_left_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[3] = chanx_left_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[4] = chanx_left_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[5] = chanx_left_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[6] = chanx_left_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[7] = chanx_left_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[8] = chanx_left_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[9] = chanx_left_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[10] = chanx_left_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[11] = chanx_left_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[12] = chanx_left_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[13] = chanx_left_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[14] = chanx_left_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[15] = chanx_left_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[16] = chanx_left_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[17] = chanx_left_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[18] = chanx_left_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[19] = chanx_left_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[20] = chanx_left_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[21] = chanx_left_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[22] = chanx_left_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[23] = chanx_left_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[24] = chanx_left_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[25] = chanx_left_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[26] = chanx_left_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[27] = chanx_left_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[28] = chanx_left_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[29] = chanx_left_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[30] = chanx_left_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[31] = chanx_left_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[32] = chanx_left_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[33] = chanx_left_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[34] = chanx_left_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[35] = chanx_left_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[36] = chanx_left_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[37] = chanx_left_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[38] = chanx_left_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[39] = chanx_left_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[40] = chanx_left_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[41] = chanx_left_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[42] = chanx_left_in[42];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[43] = chanx_left_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[44] = chanx_left_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[45] = chanx_left_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[46] = chanx_left_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[47] = chanx_left_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[48] = chanx_left_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[49] = chanx_left_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[50] = chanx_left_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[51] = chanx_left_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[52] = chanx_left_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[53] = chanx_left_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[54] = chanx_left_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[55] = chanx_left_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[56] = chanx_left_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[57] = chanx_left_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[58] = chanx_left_in[58];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[59] = chanx_left_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[60] = chanx_left_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[61] = chanx_left_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[62] = chanx_left_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[63] = chanx_left_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[64] = chanx_left_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[65] = chanx_left_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[66] = chanx_left_in[66];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[67] = chanx_left_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[68] = chanx_left_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[69] = chanx_left_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[70] = chanx_left_in[70];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[71] = chanx_left_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[72] = chanx_left_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[73] = chanx_left_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[74] = chanx_left_in[74];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[75] = chanx_left_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[76] = chanx_left_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[77] = chanx_left_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[78] = chanx_left_in[78];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[79] = chanx_left_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[0] = chanx_right_in[0];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[1] = chanx_right_in[1];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[2] = chanx_right_in[2];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[3] = chanx_right_in[3];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[4] = chanx_right_in[4];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[5] = chanx_right_in[5];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[6] = chanx_right_in[6];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[7] = chanx_right_in[7];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[8] = chanx_right_in[8];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[9] = chanx_right_in[9];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[10] = chanx_right_in[10];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[11] = chanx_right_in[11];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[12] = chanx_right_in[12];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[13] = chanx_right_in[13];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[14] = chanx_right_in[14];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[15] = chanx_right_in[15];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[16] = chanx_right_in[16];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[17] = chanx_right_in[17];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[18] = chanx_right_in[18];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[19] = chanx_right_in[19];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[20] = chanx_right_in[20];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[21] = chanx_right_in[21];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[22] = chanx_right_in[22];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[23] = chanx_right_in[23];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[24] = chanx_right_in[24];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[25] = chanx_right_in[25];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[26] = chanx_right_in[26];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[27] = chanx_right_in[27];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[28] = chanx_right_in[28];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[29] = chanx_right_in[29];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[30] = chanx_right_in[30];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[31] = chanx_right_in[31];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[32] = chanx_right_in[32];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[33] = chanx_right_in[33];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[34] = chanx_right_in[34];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[35] = chanx_right_in[35];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[36] = chanx_right_in[36];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[37] = chanx_right_in[37];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[38] = chanx_right_in[38];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[39] = chanx_right_in[39];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[40] = chanx_right_in[40];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[41] = chanx_right_in[41];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[42] = chanx_right_in[42];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[43] = chanx_right_in[43];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[44] = chanx_right_in[44];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[45] = chanx_right_in[45];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[46] = chanx_right_in[46];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[47] = chanx_right_in[47];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[48] = chanx_right_in[48];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[49] = chanx_right_in[49];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[50] = chanx_right_in[50];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[51] = chanx_right_in[51];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[52] = chanx_right_in[52];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[53] = chanx_right_in[53];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[54] = chanx_right_in[54];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[55] = chanx_right_in[55];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[56] = chanx_right_in[56];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[57] = chanx_right_in[57];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[58] = chanx_right_in[58];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[59] = chanx_right_in[59];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[60] = chanx_right_in[60];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[61] = chanx_right_in[61];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[62] = chanx_right_in[62];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[63] = chanx_right_in[63];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[64] = chanx_right_in[64];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[65] = chanx_right_in[65];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[66] = chanx_right_in[66];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[67] = chanx_right_in[67];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[68] = chanx_right_in[68];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[69] = chanx_right_in[69];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[70] = chanx_right_in[70];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[71] = chanx_right_in[71];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[72] = chanx_right_in[72];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[73] = chanx_right_in[73];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[74] = chanx_right_in[74];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[75] = chanx_right_in[75];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[76] = chanx_right_in[76];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[77] = chanx_right_in[77];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[78] = chanx_right_in[78];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out[79] = chanx_right_in[79];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size18 mux_top_ipin_0 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[16], chanx_right_in[16], chanx_left_in[24], chanx_right_in[24], chanx_left_in[32], chanx_right_in[32], chanx_left_in[40], chanx_right_in[40], chanx_left_in[48], chanx_right_in[48], chanx_left_in[56], chanx_right_in[56], chanx_left_in[64], chanx_right_in[64], chanx_left_in[72], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size18_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_0_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_1 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[17], chanx_right_in[17], chanx_left_in[25], chanx_right_in[25], chanx_left_in[33], chanx_right_in[33], chanx_left_in[41], chanx_right_in[41], chanx_left_in[49], chanx_right_in[49], chanx_left_in[57], chanx_right_in[57], chanx_left_in[65], chanx_right_in[65], chanx_left_in[73], chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_size18_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_1_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_2 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[18], chanx_right_in[18], chanx_left_in[26], chanx_right_in[26], chanx_left_in[34], chanx_right_in[34], chanx_left_in[42], chanx_right_in[42], chanx_left_in[50], chanx_right_in[50], chanx_left_in[58], chanx_right_in[58], chanx_left_in[66], chanx_right_in[66], chanx_left_in[74], chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_size18_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_2_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_3 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[19], chanx_right_in[19], chanx_left_in[27], chanx_right_in[27], chanx_left_in[35], chanx_right_in[35], chanx_left_in[43], chanx_right_in[43], chanx_left_in[51], chanx_right_in[51], chanx_left_in[59], chanx_right_in[59], chanx_left_in[67], chanx_right_in[67], chanx_left_in[75], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size18_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_3_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_4 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[20], chanx_right_in[20], chanx_left_in[28], chanx_right_in[28], chanx_left_in[36], chanx_right_in[36], chanx_left_in[44], chanx_right_in[44], chanx_left_in[52], chanx_right_in[52], chanx_left_in[60], chanx_right_in[60], chanx_left_in[68], chanx_right_in[68], chanx_left_in[76], chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_size18_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_4_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_5 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[21], chanx_right_in[21], chanx_left_in[29], chanx_right_in[29], chanx_left_in[37], chanx_right_in[37], chanx_left_in[45], chanx_right_in[45], chanx_left_in[53], chanx_right_in[53], chanx_left_in[61], chanx_right_in[61], chanx_left_in[69], chanx_right_in[69], chanx_left_in[77], chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_size18_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_5_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_6 (
		.in({chanx_left_in[6], chanx_right_in[6], chanx_left_in[22], chanx_right_in[22], chanx_left_in[30], chanx_right_in[30], chanx_left_in[38], chanx_right_in[38], chanx_left_in[46], chanx_right_in[46], chanx_left_in[54], chanx_right_in[54], chanx_left_in[62], chanx_right_in[62], chanx_left_in[70], chanx_right_in[70], chanx_left_in[78], chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_size18_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_6_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_7 (
		.in({chanx_left_in[7], chanx_right_in[7], chanx_left_in[23], chanx_right_in[23], chanx_left_in[31], chanx_right_in[31], chanx_left_in[39], chanx_right_in[39], chanx_left_in[47], chanx_right_in[47], chanx_left_in[55], chanx_right_in[55], chanx_left_in[63], chanx_right_in[63], chanx_left_in[71], chanx_right_in[71], chanx_left_in[79], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size18_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_7_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_8 (
		.in({chanx_left_in[8], chanx_right_in[8], chanx_left_in[16], chanx_right_in[16], chanx_left_in[24], chanx_right_in[24], chanx_left_in[32], chanx_right_in[32], chanx_left_in[40], chanx_right_in[40], chanx_left_in[48], chanx_right_in[48], chanx_left_in[56], chanx_right_in[56], chanx_left_in[64], chanx_right_in[64], chanx_left_in[72], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size18_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_8_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_9 (
		.in({chanx_left_in[9], chanx_right_in[9], chanx_left_in[17], chanx_right_in[17], chanx_left_in[25], chanx_right_in[25], chanx_left_in[33], chanx_right_in[33], chanx_left_in[41], chanx_right_in[41], chanx_left_in[49], chanx_right_in[49], chanx_left_in[57], chanx_right_in[57], chanx_left_in[65], chanx_right_in[65], chanx_left_in[73], chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_size18_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_9_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_10 (
		.in({chanx_left_in[10], chanx_right_in[10], chanx_left_in[18], chanx_right_in[18], chanx_left_in[26], chanx_right_in[26], chanx_left_in[34], chanx_right_in[34], chanx_left_in[42], chanx_right_in[42], chanx_left_in[50], chanx_right_in[50], chanx_left_in[58], chanx_right_in[58], chanx_left_in[66], chanx_right_in[66], chanx_left_in[74], chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_size18_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_10_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_11 (
		.in({chanx_left_in[11], chanx_right_in[11], chanx_left_in[19], chanx_right_in[19], chanx_left_in[27], chanx_right_in[27], chanx_left_in[35], chanx_right_in[35], chanx_left_in[43], chanx_right_in[43], chanx_left_in[51], chanx_right_in[51], chanx_left_in[59], chanx_right_in[59], chanx_left_in[67], chanx_right_in[67], chanx_left_in[75], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size18_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_11_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_12 (
		.in({chanx_left_in[12], chanx_right_in[12], chanx_left_in[20], chanx_right_in[20], chanx_left_in[28], chanx_right_in[28], chanx_left_in[36], chanx_right_in[36], chanx_left_in[44], chanx_right_in[44], chanx_left_in[52], chanx_right_in[52], chanx_left_in[60], chanx_right_in[60], chanx_left_in[68], chanx_right_in[68], chanx_left_in[76], chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_size18_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_12_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_13 (
		.in({chanx_left_in[13], chanx_right_in[13], chanx_left_in[21], chanx_right_in[21], chanx_left_in[29], chanx_right_in[29], chanx_left_in[37], chanx_right_in[37], chanx_left_in[45], chanx_right_in[45], chanx_left_in[53], chanx_right_in[53], chanx_left_in[61], chanx_right_in[61], chanx_left_in[69], chanx_right_in[69], chanx_left_in[77], chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_size18_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_13_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_14 (
		.in({chanx_left_in[14], chanx_right_in[14], chanx_left_in[22], chanx_right_in[22], chanx_left_in[30], chanx_right_in[30], chanx_left_in[38], chanx_right_in[38], chanx_left_in[46], chanx_right_in[46], chanx_left_in[54], chanx_right_in[54], chanx_left_in[62], chanx_right_in[62], chanx_left_in[70], chanx_right_in[70], chanx_left_in[78], chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_size18_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_14_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_15 (
		.in({chanx_left_in[15], chanx_right_in[15], chanx_left_in[23], chanx_right_in[23], chanx_left_in[31], chanx_right_in[31], chanx_left_in[39], chanx_right_in[39], chanx_left_in[47], chanx_right_in[47], chanx_left_in[55], chanx_right_in[55], chanx_left_in[63], chanx_right_in[63], chanx_left_in[71], chanx_right_in[71], chanx_left_in[79], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size18_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_15_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_16 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[16], chanx_right_in[16], chanx_left_in[24], chanx_right_in[24], chanx_left_in[32], chanx_right_in[32], chanx_left_in[40], chanx_right_in[40], chanx_left_in[48], chanx_right_in[48], chanx_left_in[56], chanx_right_in[56], chanx_left_in[64], chanx_right_in[64], chanx_left_in[72], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size18_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_16_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_17 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[17], chanx_right_in[17], chanx_left_in[25], chanx_right_in[25], chanx_left_in[33], chanx_right_in[33], chanx_left_in[41], chanx_right_in[41], chanx_left_in[49], chanx_right_in[49], chanx_left_in[57], chanx_right_in[57], chanx_left_in[65], chanx_right_in[65], chanx_left_in[73], chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_size18_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_17_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_18 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[18], chanx_right_in[18], chanx_left_in[26], chanx_right_in[26], chanx_left_in[34], chanx_right_in[34], chanx_left_in[42], chanx_right_in[42], chanx_left_in[50], chanx_right_in[50], chanx_left_in[58], chanx_right_in[58], chanx_left_in[66], chanx_right_in[66], chanx_left_in[74], chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_size18_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_18_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_19 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[19], chanx_right_in[19], chanx_left_in[27], chanx_right_in[27], chanx_left_in[35], chanx_right_in[35], chanx_left_in[43], chanx_right_in[43], chanx_left_in[51], chanx_right_in[51], chanx_left_in[59], chanx_right_in[59], chanx_left_in[67], chanx_right_in[67], chanx_left_in[75], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size18_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_19_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_20 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[20], chanx_right_in[20], chanx_left_in[28], chanx_right_in[28], chanx_left_in[36], chanx_right_in[36], chanx_left_in[44], chanx_right_in[44], chanx_left_in[52], chanx_right_in[52], chanx_left_in[60], chanx_right_in[60], chanx_left_in[68], chanx_right_in[68], chanx_left_in[76], chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_size18_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_20_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_20__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_21 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[21], chanx_right_in[21], chanx_left_in[29], chanx_right_in[29], chanx_left_in[37], chanx_right_in[37], chanx_left_in[45], chanx_right_in[45], chanx_left_in[53], chanx_right_in[53], chanx_left_in[61], chanx_right_in[61], chanx_left_in[69], chanx_right_in[69], chanx_left_in[77], chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_size18_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_21_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_21__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_22 (
		.in({chanx_left_in[6], chanx_right_in[6], chanx_left_in[22], chanx_right_in[22], chanx_left_in[30], chanx_right_in[30], chanx_left_in[38], chanx_right_in[38], chanx_left_in[46], chanx_right_in[46], chanx_left_in[54], chanx_right_in[54], chanx_left_in[62], chanx_right_in[62], chanx_left_in[70], chanx_right_in[70], chanx_left_in[78], chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_size18_22_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_22_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_22__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_23 (
		.in({chanx_left_in[7], chanx_right_in[7], chanx_left_in[23], chanx_right_in[23], chanx_left_in[31], chanx_right_in[31], chanx_left_in[39], chanx_right_in[39], chanx_left_in[47], chanx_right_in[47], chanx_left_in[55], chanx_right_in[55], chanx_left_in[63], chanx_right_in[63], chanx_left_in[71], chanx_right_in[71], chanx_left_in[79], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size18_23_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_23_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_23__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_24 (
		.in({chanx_left_in[8], chanx_right_in[8], chanx_left_in[16], chanx_right_in[16], chanx_left_in[24], chanx_right_in[24], chanx_left_in[32], chanx_right_in[32], chanx_left_in[40], chanx_right_in[40], chanx_left_in[48], chanx_right_in[48], chanx_left_in[56], chanx_right_in[56], chanx_left_in[64], chanx_right_in[64], chanx_left_in[72], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size18_24_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_24_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_24__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_25 (
		.in({chanx_left_in[9], chanx_right_in[9], chanx_left_in[17], chanx_right_in[17], chanx_left_in[25], chanx_right_in[25], chanx_left_in[33], chanx_right_in[33], chanx_left_in[41], chanx_right_in[41], chanx_left_in[49], chanx_right_in[49], chanx_left_in[57], chanx_right_in[57], chanx_left_in[65], chanx_right_in[65], chanx_left_in[73], chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_size18_25_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_25_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_25__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_26 (
		.in({chanx_left_in[10], chanx_right_in[10], chanx_left_in[18], chanx_right_in[18], chanx_left_in[26], chanx_right_in[26], chanx_left_in[34], chanx_right_in[34], chanx_left_in[42], chanx_right_in[42], chanx_left_in[50], chanx_right_in[50], chanx_left_in[58], chanx_right_in[58], chanx_left_in[66], chanx_right_in[66], chanx_left_in[74], chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_size18_26_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_26_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_26__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_27 (
		.in({chanx_left_in[11], chanx_right_in[11], chanx_left_in[19], chanx_right_in[19], chanx_left_in[27], chanx_right_in[27], chanx_left_in[35], chanx_right_in[35], chanx_left_in[43], chanx_right_in[43], chanx_left_in[51], chanx_right_in[51], chanx_left_in[59], chanx_right_in[59], chanx_left_in[67], chanx_right_in[67], chanx_left_in[75], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size18_27_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_27_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_27__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_28 (
		.in({chanx_left_in[12], chanx_right_in[12], chanx_left_in[20], chanx_right_in[20], chanx_left_in[28], chanx_right_in[28], chanx_left_in[36], chanx_right_in[36], chanx_left_in[44], chanx_right_in[44], chanx_left_in[52], chanx_right_in[52], chanx_left_in[60], chanx_right_in[60], chanx_left_in[68], chanx_right_in[68], chanx_left_in[76], chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_size18_28_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_28_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_28__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_29 (
		.in({chanx_left_in[13], chanx_right_in[13], chanx_left_in[21], chanx_right_in[21], chanx_left_in[29], chanx_right_in[29], chanx_left_in[37], chanx_right_in[37], chanx_left_in[45], chanx_right_in[45], chanx_left_in[53], chanx_right_in[53], chanx_left_in[61], chanx_right_in[61], chanx_left_in[69], chanx_right_in[69], chanx_left_in[77], chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_size18_29_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_29_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_29__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_30 (
		.in({chanx_left_in[14], chanx_right_in[14], chanx_left_in[22], chanx_right_in[22], chanx_left_in[30], chanx_right_in[30], chanx_left_in[38], chanx_right_in[38], chanx_left_in[46], chanx_right_in[46], chanx_left_in[54], chanx_right_in[54], chanx_left_in[62], chanx_right_in[62], chanx_left_in[70], chanx_right_in[70], chanx_left_in[78], chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_size18_30_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_30_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_30__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_31 (
		.in({chanx_left_in[15], chanx_right_in[15], chanx_left_in[23], chanx_right_in[23], chanx_left_in[31], chanx_right_in[31], chanx_left_in[39], chanx_right_in[39], chanx_left_in[47], chanx_right_in[47], chanx_left_in[55], chanx_right_in[55], chanx_left_in[63], chanx_right_in[63], chanx_left_in[71], chanx_right_in[71], chanx_left_in[79], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size18_31_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_31_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_31__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_32 (
		.in({chanx_left_in[0], chanx_right_in[0], chanx_left_in[16], chanx_right_in[16], chanx_left_in[24], chanx_right_in[24], chanx_left_in[32], chanx_right_in[32], chanx_left_in[40], chanx_right_in[40], chanx_left_in[48], chanx_right_in[48], chanx_left_in[56], chanx_right_in[56], chanx_left_in[64], chanx_right_in[64], chanx_left_in[72], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size18_32_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_32_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_32__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_33 (
		.in({chanx_left_in[1], chanx_right_in[1], chanx_left_in[17], chanx_right_in[17], chanx_left_in[25], chanx_right_in[25], chanx_left_in[33], chanx_right_in[33], chanx_left_in[41], chanx_right_in[41], chanx_left_in[49], chanx_right_in[49], chanx_left_in[57], chanx_right_in[57], chanx_left_in[65], chanx_right_in[65], chanx_left_in[73], chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_size18_33_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_33_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_33__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_34 (
		.in({chanx_left_in[2], chanx_right_in[2], chanx_left_in[18], chanx_right_in[18], chanx_left_in[26], chanx_right_in[26], chanx_left_in[34], chanx_right_in[34], chanx_left_in[42], chanx_right_in[42], chanx_left_in[50], chanx_right_in[50], chanx_left_in[58], chanx_right_in[58], chanx_left_in[66], chanx_right_in[66], chanx_left_in[74], chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_size18_34_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_34_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_34__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_35 (
		.in({chanx_left_in[3], chanx_right_in[3], chanx_left_in[19], chanx_right_in[19], chanx_left_in[27], chanx_right_in[27], chanx_left_in[35], chanx_right_in[35], chanx_left_in[43], chanx_right_in[43], chanx_left_in[51], chanx_right_in[51], chanx_left_in[59], chanx_right_in[59], chanx_left_in[67], chanx_right_in[67], chanx_left_in[75], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size18_35_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_35_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_35__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_36 (
		.in({chanx_left_in[4], chanx_right_in[4], chanx_left_in[20], chanx_right_in[20], chanx_left_in[28], chanx_right_in[28], chanx_left_in[36], chanx_right_in[36], chanx_left_in[44], chanx_right_in[44], chanx_left_in[52], chanx_right_in[52], chanx_left_in[60], chanx_right_in[60], chanx_left_in[68], chanx_right_in[68], chanx_left_in[76], chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_size18_36_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_36_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_36__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_37 (
		.in({chanx_left_in[5], chanx_right_in[5], chanx_left_in[21], chanx_right_in[21], chanx_left_in[29], chanx_right_in[29], chanx_left_in[37], chanx_right_in[37], chanx_left_in[45], chanx_right_in[45], chanx_left_in[53], chanx_right_in[53], chanx_left_in[61], chanx_right_in[61], chanx_left_in[69], chanx_right_in[69], chanx_left_in[77], chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_size18_37_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_37_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_37__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_38 (
		.in({chanx_left_in[6], chanx_right_in[6], chanx_left_in[22], chanx_right_in[22], chanx_left_in[30], chanx_right_in[30], chanx_left_in[38], chanx_right_in[38], chanx_left_in[46], chanx_right_in[46], chanx_left_in[54], chanx_right_in[54], chanx_left_in[62], chanx_right_in[62], chanx_left_in[70], chanx_right_in[70], chanx_left_in[78], chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_size18_38_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_38_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_38__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_39 (
		.in({chanx_left_in[7], chanx_right_in[7], chanx_left_in[23], chanx_right_in[23], chanx_left_in[31], chanx_right_in[31], chanx_left_in[39], chanx_right_in[39], chanx_left_in[47], chanx_right_in[47], chanx_left_in[55], chanx_right_in[55], chanx_left_in[63], chanx_right_in[63], chanx_left_in[71], chanx_right_in[71], chanx_left_in[79], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size18_39_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_39_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_39__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_40 (
		.in({chanx_left_in[8], chanx_right_in[8], chanx_left_in[16], chanx_right_in[16], chanx_left_in[24], chanx_right_in[24], chanx_left_in[32], chanx_right_in[32], chanx_left_in[40], chanx_right_in[40], chanx_left_in[48], chanx_right_in[48], chanx_left_in[56], chanx_right_in[56], chanx_left_in[64], chanx_right_in[64], chanx_left_in[72], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size18_40_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_40_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_40__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_41 (
		.in({chanx_left_in[9], chanx_right_in[9], chanx_left_in[17], chanx_right_in[17], chanx_left_in[25], chanx_right_in[25], chanx_left_in[33], chanx_right_in[33], chanx_left_in[41], chanx_right_in[41], chanx_left_in[49], chanx_right_in[49], chanx_left_in[57], chanx_right_in[57], chanx_left_in[65], chanx_right_in[65], chanx_left_in[73], chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_size18_41_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_41_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_41__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_42 (
		.in({chanx_left_in[10], chanx_right_in[10], chanx_left_in[18], chanx_right_in[18], chanx_left_in[26], chanx_right_in[26], chanx_left_in[34], chanx_right_in[34], chanx_left_in[42], chanx_right_in[42], chanx_left_in[50], chanx_right_in[50], chanx_left_in[58], chanx_right_in[58], chanx_left_in[66], chanx_right_in[66], chanx_left_in[74], chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_size18_42_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_42_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_42__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_43 (
		.in({chanx_left_in[11], chanx_right_in[11], chanx_left_in[19], chanx_right_in[19], chanx_left_in[27], chanx_right_in[27], chanx_left_in[35], chanx_right_in[35], chanx_left_in[43], chanx_right_in[43], chanx_left_in[51], chanx_right_in[51], chanx_left_in[59], chanx_right_in[59], chanx_left_in[67], chanx_right_in[67], chanx_left_in[75], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size18_43_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_43_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_43__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_44 (
		.in({chanx_left_in[12], chanx_right_in[12], chanx_left_in[20], chanx_right_in[20], chanx_left_in[28], chanx_right_in[28], chanx_left_in[36], chanx_right_in[36], chanx_left_in[44], chanx_right_in[44], chanx_left_in[52], chanx_right_in[52], chanx_left_in[60], chanx_right_in[60], chanx_left_in[68], chanx_right_in[68], chanx_left_in[76], chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_size18_44_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_44_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_44__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_45 (
		.in({chanx_left_in[13], chanx_right_in[13], chanx_left_in[21], chanx_right_in[21], chanx_left_in[29], chanx_right_in[29], chanx_left_in[37], chanx_right_in[37], chanx_left_in[45], chanx_right_in[45], chanx_left_in[53], chanx_right_in[53], chanx_left_in[61], chanx_right_in[61], chanx_left_in[69], chanx_right_in[69], chanx_left_in[77], chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_size18_45_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_45_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_45__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_46 (
		.in({chanx_left_in[14], chanx_right_in[14], chanx_left_in[22], chanx_right_in[22], chanx_left_in[30], chanx_right_in[30], chanx_left_in[38], chanx_right_in[38], chanx_left_in[46], chanx_right_in[46], chanx_left_in[54], chanx_right_in[54], chanx_left_in[62], chanx_right_in[62], chanx_left_in[70], chanx_right_in[70], chanx_left_in[78], chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_size18_46_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_46_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_46__pin_f2a_i_0_));

	mux_tree_tapbuf_size18 mux_top_ipin_47 (
		.in({chanx_left_in[15], chanx_right_in[15], chanx_left_in[23], chanx_right_in[23], chanx_left_in[31], chanx_right_in[31], chanx_left_in[39], chanx_right_in[39], chanx_left_in[47], chanx_right_in[47], chanx_left_in[55], chanx_right_in[55], chanx_left_in[63], chanx_right_in[63], chanx_left_in[71], chanx_right_in[71], chanx_left_in[79], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size18_47_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_47_sram_inv[0:4]),
		.out(bottom_grid_top_width_0_height_0_subtile_47__pin_f2a_i_0_));

	mux_tree_tapbuf_size18_mem mem_top_ipin_0 (
		.bl(bl[0:4]),
		.wl({wl[0], wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_size18_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_0_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_1 (
		.bl(bl[5:9]),
		.wl({wl[0], wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_size18_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_1_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_2 (
		.bl(bl[10:14]),
		.wl({wl[0], wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_size18_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_2_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_3 (
		.bl({bl[15], bl[0:3]}),
		.wl({wl[0:1], wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_size18_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_3_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_4 (
		.bl(bl[4:8]),
		.wl({wl[1], wl[1], wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_size18_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_4_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_5 (
		.bl(bl[9:13]),
		.wl({wl[1], wl[1], wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_size18_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_5_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_6 (
		.bl({bl[14:15], bl[0:2]}),
		.wl({wl[1], wl[1:2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_size18_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_6_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_7 (
		.bl(bl[3:7]),
		.wl({wl[2], wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_size18_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_7_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_8 (
		.bl(bl[8:12]),
		.wl({wl[2], wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_size18_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_8_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_9 (
		.bl({bl[13:15], bl[0:1]}),
		.wl({wl[2], wl[2], wl[2:3], wl[3]}),
		.mem_out(mux_tree_tapbuf_size18_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_9_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_10 (
		.bl(bl[2:6]),
		.wl({wl[3], wl[3], wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_size18_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_10_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_11 (
		.bl(bl[7:11]),
		.wl({wl[3], wl[3], wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_size18_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_11_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_12 (
		.bl({bl[12:15], bl[0]}),
		.wl({wl[3], wl[3], wl[3], wl[3:4]}),
		.mem_out(mux_tree_tapbuf_size18_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_12_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_13 (
		.bl(bl[1:5]),
		.wl({wl[4], wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_size18_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_13_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_14 (
		.bl(bl[6:10]),
		.wl({wl[4], wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_size18_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_14_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_15 (
		.bl(bl[11:15]),
		.wl({wl[4], wl[4], wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_size18_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_15_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_16 (
		.bl(bl[0:4]),
		.wl({wl[5], wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_size18_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_16_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_17 (
		.bl(bl[5:9]),
		.wl({wl[5], wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_size18_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_17_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_18 (
		.bl(bl[10:14]),
		.wl({wl[5], wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_size18_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_18_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_19 (
		.bl({bl[15], bl[0:3]}),
		.wl({wl[5:6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_size18_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_19_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_20 (
		.bl(bl[4:8]),
		.wl({wl[6], wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_size18_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_20_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_21 (
		.bl(bl[9:13]),
		.wl({wl[6], wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_size18_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_21_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_22 (
		.bl({bl[14:15], bl[0:2]}),
		.wl({wl[6], wl[6:7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_size18_22_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_22_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_23 (
		.bl(bl[3:7]),
		.wl({wl[7], wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_size18_23_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_23_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_24 (
		.bl(bl[8:12]),
		.wl({wl[7], wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_size18_24_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_24_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_25 (
		.bl({bl[13:15], bl[0:1]}),
		.wl({wl[7], wl[7], wl[7:8], wl[8]}),
		.mem_out(mux_tree_tapbuf_size18_25_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_25_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_26 (
		.bl(bl[2:6]),
		.wl({wl[8], wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_size18_26_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_26_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_27 (
		.bl(bl[7:11]),
		.wl({wl[8], wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_size18_27_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_27_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_28 (
		.bl({bl[12:15], bl[0]}),
		.wl({wl[8], wl[8], wl[8], wl[8:9]}),
		.mem_out(mux_tree_tapbuf_size18_28_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_28_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_29 (
		.bl(bl[1:5]),
		.wl({wl[9], wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_size18_29_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_29_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_30 (
		.bl(bl[6:10]),
		.wl({wl[9], wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_size18_30_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_30_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_31 (
		.bl(bl[11:15]),
		.wl({wl[9], wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_size18_31_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_31_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_32 (
		.bl(bl[0:4]),
		.wl({wl[10], wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_size18_32_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_32_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_33 (
		.bl(bl[5:9]),
		.wl({wl[10], wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_size18_33_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_33_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_34 (
		.bl(bl[10:14]),
		.wl({wl[10], wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_size18_34_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_34_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_35 (
		.bl({bl[15], bl[0:3]}),
		.wl({wl[10:11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_size18_35_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_35_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_36 (
		.bl(bl[4:8]),
		.wl({wl[11], wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_size18_36_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_36_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_37 (
		.bl(bl[9:13]),
		.wl({wl[11], wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_size18_37_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_37_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_38 (
		.bl({bl[14:15], bl[0:2]}),
		.wl({wl[11], wl[11:12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_size18_38_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_38_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_39 (
		.bl(bl[3:7]),
		.wl({wl[12], wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_size18_39_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_39_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_40 (
		.bl(bl[8:12]),
		.wl({wl[12], wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_size18_40_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_40_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_41 (
		.bl({bl[13:15], bl[0:1]}),
		.wl({wl[12], wl[12], wl[12:13], wl[13]}),
		.mem_out(mux_tree_tapbuf_size18_41_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_41_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_42 (
		.bl(bl[2:6]),
		.wl({wl[13], wl[13], wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_size18_42_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_42_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_43 (
		.bl(bl[7:11]),
		.wl({wl[13], wl[13], wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_size18_43_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_43_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_44 (
		.bl({bl[12:15], bl[0]}),
		.wl({wl[13], wl[13], wl[13], wl[13:14]}),
		.mem_out(mux_tree_tapbuf_size18_44_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_44_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_45 (
		.bl(bl[1:5]),
		.wl({wl[14], wl[14], wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_size18_45_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_45_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_46 (
		.bl(bl[6:10]),
		.wl({wl[14], wl[14], wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_size18_46_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_46_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_ipin_47 (
		.bl(bl[11:15]),
		.wl({wl[14], wl[14], wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_size18_47_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_47_sram_inv[0:4]));

endmodule
// ----- END Verilog module for cbx_1__1_ -----

//----- Default net type -----
`default_nettype none




