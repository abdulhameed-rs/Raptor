//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][1]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_1__1_ -----
module sb_1__1_(chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                chanx_right_in,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_,
                chany_bottom_in,
                bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                chanx_left_in,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_,
                bl,
                wl,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out);
//----- INPUT PORTS -----
input [0:79] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:79] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:79] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:79] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:21] bl;
//----- INPUT PORTS -----
input [0:21] wl;
//----- OUTPUT PORTS -----
output [0:79] chany_top_out;
//----- OUTPUT PORTS -----
output [0:79] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:79] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:79] chanx_left_out;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_L1SB_size11_0_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size11_1_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size11_2_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size11_3_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size11_4_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size11_5_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size11_6_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size11_7_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_0_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_10_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_11_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_12_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_13_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_14_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_15_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_16_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_16_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_17_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_17_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_18_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_18_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_19_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_19_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_1_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_20_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_20_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_21_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_21_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_22_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_22_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_23_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_23_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_2_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_3_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_4_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_5_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_6_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_7_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_8_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size12_9_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size12_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_2_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_3_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_4_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_5_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_6_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_7_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_0_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_10_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_11_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_12_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_13_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_14_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_15_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_16_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_16_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_17_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_17_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_18_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_18_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_19_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_19_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_1_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_20_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_20_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_21_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_21_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_22_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_22_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_23_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_23_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_2_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_3_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_4_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_5_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_6_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_7_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_8_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_9_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_14_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_15_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_14_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_15_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L1SB_size9 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, chanx_right_in[1], chanx_right_in[16], chanx_right_in[58], chany_bottom_in[16], chany_bottom_in[58], chanx_left_in[0], chanx_left_in[16], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L1SB_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_0_sram_inv[0:3]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, chanx_right_in[2], chanx_right_in[17], chanx_right_in[60], chany_bottom_in[17], chany_bottom_in[60], chanx_left_in[17], chanx_left_in[60], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L1SB_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_1_sram_inv[0:3]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, chanx_right_in[3], chanx_right_in[18], chanx_right_in[61], chany_bottom_in[18], chany_bottom_in[61], chanx_left_in[18], chanx_left_in[61], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L1SB_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_2_sram_inv[0:3]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, chanx_right_in[4], chanx_right_in[20], chanx_right_in[62], chany_bottom_in[20], chany_bottom_in[62], chanx_left_in[20], chanx_left_in[62], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L1SB_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_3_sram_inv[0:3]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_right_in[5], chanx_right_in[21], chanx_right_in[64], chany_bottom_in[21], chany_bottom_in[64], chanx_left_in[21], chanx_left_in[64], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L1SB_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_4_sram_inv[0:3]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_right_in[6], chanx_right_in[22], chanx_right_in[65], chany_bottom_in[22], chany_bottom_in[65], chanx_left_in[22], chanx_left_in[63], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L1SB_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_5_sram_inv[0:3]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_right_in[7], chanx_right_in[24], chanx_right_in[66], chany_bottom_in[24], chany_bottom_in[66], chanx_left_in[24], chanx_left_in[59], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L1SB_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_6_sram_inv[0:3]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[8], chanx_right_in[25], chanx_right_in[68], chany_bottom_in[25], chany_bottom_in[68], chanx_left_in[25], chanx_left_in[55], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L1SB_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_7_sram_inv[0:3]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_right_in[9], chanx_right_in[26], chanx_right_in[69], chany_bottom_in[26], chany_bottom_in[69], chanx_left_in[26], chanx_left_in[51], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L1SB_size9_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_8_sram_inv[0:3]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_right_in[10], chanx_right_in[28], chanx_right_in[70], chany_bottom_in[28], chany_bottom_in[70], chanx_left_in[28], chanx_left_in[47], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L1SB_size9_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_9_sram_inv[0:3]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_right_in[11], chanx_right_in[29], chanx_right_in[72], chany_bottom_in[29], chany_bottom_in[72], chanx_left_in[29], chanx_left_in[43], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size9_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_10_sram_inv[0:3]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_L1SB_size9 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_right_in[12], chanx_right_in[30], chanx_right_in[73], chany_bottom_in[30], chany_bottom_in[73], chanx_left_in[30], chanx_left_in[39], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size9_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_11_sram_inv[0:3]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_1 (
		.in({chany_top_in[16], chany_top_in[58], chanx_right_in[16], chanx_right_in[58], chanx_right_in[75], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, chanx_left_in[1], chanx_left_in[16], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L1SB_size9_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_12_sram_inv[0:3]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_3 (
		.in({chany_top_in[17], chany_top_in[60], chanx_right_in[17], chanx_right_in[60], chanx_right_in[71], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, chanx_left_in[2], chanx_left_in[17], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L1SB_size9_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_13_sram_inv[0:3]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_5 (
		.in({chany_top_in[18], chany_top_in[61], chanx_right_in[18], chanx_right_in[61], chanx_right_in[67], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, chanx_left_in[3], chanx_left_in[18], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L1SB_size9_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_14_sram_inv[0:3]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_7 (
		.in({chany_top_in[20], chany_top_in[62], chanx_right_in[20], chanx_right_in[62:63], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, chanx_left_in[4], chanx_left_in[20], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L1SB_size9_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_15_sram_inv[0:3]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_9 (
		.in({chany_top_in[21], chany_top_in[64], chanx_right_in[21], chanx_right_in[59], chanx_right_in[64], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_left_in[5], chanx_left_in[21], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L1SB_size9_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_16_sram_inv[0:3]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_11 (
		.in({chany_top_in[22], chany_top_in[65], chanx_right_in[22], chanx_right_in[55], chanx_right_in[65], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[6], chanx_left_in[22], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L1SB_size9_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_17_sram_inv[0:3]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_13 (
		.in({chany_top_in[24], chany_top_in[66], chanx_right_in[24], chanx_right_in[51], chanx_right_in[66], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[7], chanx_left_in[24], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L1SB_size9_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_18_sram_inv[0:3]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_15 (
		.in({chany_top_in[25], chany_top_in[68], chanx_right_in[25], chanx_right_in[47], chanx_right_in[68], bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[8], chanx_left_in[25], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L1SB_size9_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_19_sram_inv[0:3]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_17 (
		.in({chany_top_in[26], chany_top_in[69], chanx_right_in[26], chanx_right_in[43], chanx_right_in[69], bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[9], chanx_left_in[26], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L1SB_size9_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_20_sram_inv[0:3]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_19 (
		.in({chany_top_in[28], chany_top_in[70], chanx_right_in[28], chanx_right_in[39], chanx_right_in[70], bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[10], chanx_left_in[28], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L1SB_size9_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_21_sram_inv[0:3]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_21 (
		.in({chany_top_in[29], chany_top_in[72], chanx_right_in[29], chanx_right_in[35], chanx_right_in[72], bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[11], chanx_left_in[29], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size9_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_22_sram_inv[0:3]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_23 (
		.in({chany_top_in[30], chany_top_in[73], chanx_right_in[30:31], chanx_right_in[73], bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[12], chanx_left_in[30], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size9_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_23_sram_inv[0:3]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_0 (
		.bl(bl[0:3]),
		.wl({wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_2 (
		.bl(bl[4:7]),
		.wl({wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_4 (
		.bl(bl[8:11]),
		.wl({wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_6 (
		.bl(bl[12:15]),
		.wl({wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_8 (
		.bl(bl[16:19]),
		.wl({wl[0], wl[0], wl[0], wl[0]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_10 (
		.bl({bl[20:21], bl[0:1]}),
		.wl({wl[0], wl[0:1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_12 (
		.bl(bl[2:5]),
		.wl({wl[1], wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_14 (
		.bl(bl[6:9]),
		.wl({wl[1], wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_16 (
		.bl(bl[10:13]),
		.wl({wl[1], wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_8_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_18 (
		.bl(bl[14:17]),
		.wl({wl[1], wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_9_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_20 (
		.bl(bl[18:21]),
		.wl({wl[1], wl[1], wl[1], wl[1]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_10_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_top_track_22 (
		.bl(bl[0:3]),
		.wl({wl[2], wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_11_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_1 (
		.bl(bl[16:19]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_12_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_3 (
		.bl({bl[20:21], bl[0:1]}),
		.wl({wl[10], wl[10:11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_13_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_5 (
		.bl(bl[2:5]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_14_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_7 (
		.bl(bl[6:9]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_15_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_9 (
		.bl(bl[10:13]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_16_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_11 (
		.bl(bl[14:17]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_17_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_13 (
		.bl(bl[18:21]),
		.wl({wl[11], wl[11], wl[11], wl[11]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_18_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_15 (
		.bl(bl[0:3]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_19_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_17 (
		.bl(bl[4:7]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_20_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_19 (
		.bl(bl[8:11]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_21_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_21 (
		.bl(bl[12:15]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_22_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_23 (
		.bl(bl[16:19]),
		.wl({wl[12], wl[12], wl[12], wl[12]}),
		.mem_out(mux_tree_tapbuf_L1SB_size9_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_23_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_24 (
		.in({chanx_right_in[13], chanx_right_in[32], chanx_right_in[74], chany_bottom_in[32], chany_bottom_in[74], chanx_left_in[32], chanx_left_in[35], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L1SB_size8_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_0_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_26 (
		.in({chanx_right_in[14], chanx_right_in[33], chanx_right_in[76], chany_bottom_in[33], chany_bottom_in[76], chanx_left_in[31], chanx_left_in[33], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size8_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_1_sram_inv[0:2]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_28 (
		.in({chanx_right_in[15], chanx_right_in[34], chanx_right_in[77], chany_bottom_in[34], chany_bottom_in[77], chanx_left_in[27], chanx_left_in[34], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size8_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_2_sram_inv[0:2]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_30 (
		.in({chanx_right_in[19], chanx_right_in[36], chanx_right_in[78], chany_bottom_in[36], chany_bottom_in[78], chanx_left_in[23], chanx_left_in[36], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L1SB_size8_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_3_sram_inv[0:2]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_25 (
		.in({chany_top_in[32], chany_top_in[74], chanx_right_in[27], chanx_right_in[32], chanx_right_in[74], chanx_left_in[13], chanx_left_in[32], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L1SB_size8_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_4_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_27 (
		.in({chany_top_in[33], chany_top_in[76], chanx_right_in[23], chanx_right_in[33], chanx_right_in[76], chanx_left_in[14], chanx_left_in[33], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size8_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_5_sram_inv[0:2]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_29 (
		.in({chany_top_in[34], chany_top_in[77], chanx_right_in[19], chanx_right_in[34], chanx_right_in[77], chanx_left_in[15], chanx_left_in[34], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size8_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_6_sram_inv[0:2]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_31 (
		.in({chany_top_in[36], chany_top_in[78], chanx_right_in[15], chanx_right_in[36], chanx_right_in[78], chanx_left_in[19], chanx_left_in[36], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L1SB_size8_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_7_sram_inv[0:2]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_24 (
		.bl(bl[4:6]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_26 (
		.bl(bl[7:9]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_1_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_28 (
		.bl(bl[10:12]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_2_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_30 (
		.bl(bl[13:15]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_3_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_25 (
		.bl({bl[20:21], bl[0]}),
		.wl({wl[12], wl[12:13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_4_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_27 (
		.bl(bl[1:3]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_5_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_29 (
		.bl(bl[4:6]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_6_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_31 (
		.bl(bl[7:9]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L1SB_size8_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_right_in[23], chanx_right_in[37], chany_bottom_in[37], chanx_left_in[19], chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_right_in[27], chanx_right_in[38], chany_bottom_in[38], chanx_left_in[15], chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_right_in[31], chanx_right_in[40], chany_bottom_in[40], chanx_left_in[14], chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_right_in[35], chanx_right_in[41], chany_bottom_in[41], chanx_left_in[13], chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_right_in[48], chanx_right_in[55], chany_bottom_in[48], chanx_left_in[8], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_right_in[49], chanx_right_in[59], chany_bottom_in[49], chanx_left_in[7], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_right_in[50], chanx_right_in[63], chany_bottom_in[50], chanx_left_in[6], chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_right_in[52], chanx_right_in[67], chany_bottom_in[52], chanx_left_in[5], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_33 (
		.in({chany_top_in[37], chanx_right_in[14], chanx_right_in[37], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[23], chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_41 (
		.in({chany_top_in[38], chanx_right_in[13], chanx_right_in[38], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[27], chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_49 (
		.in({chany_top_in[40], chanx_right_in[12], chanx_right_in[40], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[31], chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_57 (
		.in({chany_top_in[41], chanx_right_in[11], chanx_right_in[41], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[35], chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size7_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_11_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_97 (
		.in({chany_top_in[48], chanx_right_in[6], chanx_right_in[48], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[48], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size7_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_12_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_105 (
		.in({chany_top_in[49], chanx_right_in[5], chanx_right_in[49], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[49], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size7_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_13_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_113 (
		.in({chany_top_in[50], chanx_right_in[4], chanx_right_in[50], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[50], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size7_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_14_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_121 (
		.in({chany_top_in[52], chanx_right_in[3], chanx_right_in[52], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[52], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size7_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_15_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_32 (
		.bl(bl[16:18]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_40 (
		.bl(bl[19:21]),
		.wl({wl[2], wl[2], wl[2]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_48 (
		.bl(bl[0:2]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_56 (
		.bl(bl[3:5]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_96 (
		.bl(bl[18:20]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_104 (
		.bl({bl[21], bl[0:1]}),
		.wl({wl[3:4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_112 (
		.bl(bl[2:4]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_120 (
		.bl(bl[5:7]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_33 (
		.bl(bl[10:12]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_41 (
		.bl(bl[13:15]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_49 (
		.bl(bl[16:18]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_57 (
		.bl(bl[19:21]),
		.wl({wl[13], wl[13], wl[13]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_97 (
		.bl(bl[12:14]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_105 (
		.bl(bl[15:17]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_113 (
		.bl(bl[18:20]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_14_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_121 (
		.bl({bl[21], bl[0:1]}),
		.wl({wl[14:15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size7_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_15_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_right_in[39], chanx_right_in[42], chany_bottom_in[42], chanx_left_in[12], chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_0_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_L4SB_size6 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_right_in[43:44], chany_bottom_in[44], chanx_left_in[11], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_1_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_L4SB_size6 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_right_in[45], chanx_right_in[47], chany_bottom_in[45], chanx_left_in[10], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_2_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_L4SB_size6 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[46], chanx_right_in[51], chany_bottom_in[46], chanx_left_in[9], chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_3_sram_inv[0:2]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_L4SB_size6 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_right_in[53], chanx_right_in[71], chany_bottom_in[53], chanx_left_in[4], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_4_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_L4SB_size6 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_right_in[54], chanx_right_in[75], chany_bottom_in[54], chanx_left_in[3], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_5_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_L4SB_size6 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_right_in[56], chanx_right_in[79], chany_bottom_in[56], chanx_left_in[2], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_6_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_L4SB_size6 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_right_in[0], chanx_right_in[57], chany_bottom_in[57], chanx_left_in[1], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_7_sram_inv[0:2]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_65 (
		.in({chany_top_in[42], chanx_right_in[10], chanx_right_in[42], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_left_in[39], chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_8_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_73 (
		.in({chany_top_in[44], chanx_right_in[9], chanx_right_in[44], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[43:44]}),
		.sram(mux_tree_tapbuf_L4SB_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_9_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_81 (
		.in({chany_top_in[45], chanx_right_in[8], chanx_right_in[45], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[45], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_10_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_89 (
		.in({chany_top_in[46], chanx_right_in[7], chanx_right_in[46], bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[46], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size6_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_11_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_129 (
		.in({chany_top_in[53], chanx_right_in[2], chanx_right_in[53], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_left_in[53], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size6_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_12_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_137 (
		.in({chany_top_in[54], chanx_right_in[1], chanx_right_in[54], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[54], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size6_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_13_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_145 (
		.in({chany_top_in[56], chanx_right_in[0], chanx_right_in[56], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[56], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size6_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_14_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_153 (
		.in({chany_top_in[57], chanx_right_in[57], chanx_right_in[79], bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[0], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size6_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_15_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_L4SB_size6_mem mem_top_track_64 (
		.bl(bl[6:8]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_top_track_72 (
		.bl(bl[9:11]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_top_track_80 (
		.bl(bl[12:14]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_top_track_88 (
		.bl(bl[15:17]),
		.wl({wl[3], wl[3], wl[3]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_top_track_128 (
		.bl(bl[8:10]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_top_track_136 (
		.bl(bl[11:13]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_top_track_144 (
		.bl(bl[14:16]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_top_track_152 (
		.bl(bl[17:19]),
		.wl({wl[4], wl[4], wl[4]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_65 (
		.bl(bl[0:2]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_73 (
		.bl(bl[3:5]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_81 (
		.bl(bl[6:8]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_89 (
		.bl(bl[9:11]),
		.wl({wl[14], wl[14], wl[14]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_129 (
		.bl(bl[2:4]),
		.wl({wl[15], wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_137 (
		.bl(bl[5:7]),
		.wl({wl[15], wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_145 (
		.bl(bl[8:10]),
		.wl({wl[15], wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_14_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_153 (
		.bl(bl[11:13]),
		.wl({wl[15], wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L4SB_size6_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_15_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_0 (
		.in({chany_top_in[16], chany_top_in[58], chany_top_in[79], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, chany_bottom_in[16], chany_bottom_in[58], chany_bottom_in[75], chanx_left_in[16], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L1SB_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[17], chany_top_in[60], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, chany_bottom_in[17], chany_bottom_in[60], chany_bottom_in[71], chanx_left_in[17], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L1SB_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_1_sram_inv[0:3]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[18], chany_top_in[61], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, chany_bottom_in[18], chany_bottom_in[61], chany_bottom_in[67], chanx_left_in[18], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L1SB_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_2_sram_inv[0:3]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[20], chany_top_in[62], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, chany_bottom_in[20], chany_bottom_in[62:63], chanx_left_in[20], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L1SB_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_3_sram_inv[0:3]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_8 (
		.in({chany_top_in[3], chany_top_in[21], chany_top_in[64], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, chany_bottom_in[21], chany_bottom_in[59], chany_bottom_in[64], chanx_left_in[21], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L1SB_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_4_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_10 (
		.in({chany_top_in[4], chany_top_in[22], chany_top_in[65], right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, chany_bottom_in[22], chany_bottom_in[55], chany_bottom_in[65], chanx_left_in[22], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L1SB_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_5_sram_inv[0:3]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_12 (
		.in({chany_top_in[5], chany_top_in[24], chany_top_in[66], right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, chany_bottom_in[24], chany_bottom_in[51], chany_bottom_in[66], chanx_left_in[24], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L1SB_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_6_sram_inv[0:3]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_14 (
		.in({chany_top_in[6], chany_top_in[25], chany_top_in[68], right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, chany_bottom_in[25], chany_bottom_in[47], chany_bottom_in[68], chanx_left_in[25], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L1SB_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_7_sram_inv[0:3]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_16 (
		.in({chany_top_in[7], chany_top_in[26], chany_top_in[69], right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, chany_bottom_in[26], chany_bottom_in[43], chany_bottom_in[69], chanx_left_in[26], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L1SB_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_8_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_18 (
		.in({chany_top_in[8], chany_top_in[28], chany_top_in[70], right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, chany_bottom_in[28], chany_bottom_in[39], chany_bottom_in[70], chanx_left_in[28], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L1SB_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_9_sram_inv[0:3]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_20 (
		.in({chany_top_in[9], chany_top_in[29], chany_top_in[72], right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_, chany_bottom_in[29], chany_bottom_in[35], chany_bottom_in[72], chanx_left_in[29], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_10_sram_inv[0:3]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_L1SB_size12 mux_right_track_22 (
		.in({chany_top_in[10], chany_top_in[30], chany_top_in[73], right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_, chany_bottom_in[30:31], chany_bottom_in[73], chanx_left_in[30], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_11_sram_inv[0:3]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[16], chany_top_in[58], chanx_right_in[16], chanx_right_in[58], chany_bottom_in[16], chany_bottom_in[58], chany_bottom_in[79], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_12_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_3 (
		.in({chany_top_in[17], chany_top_in[60], chany_top_in[79], chanx_right_in[17], chanx_right_in[60], chany_bottom_in[0], chany_bottom_in[17], chany_bottom_in[60], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_13_sram_inv[0:3]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_5 (
		.in({chany_top_in[18], chany_top_in[61], chany_top_in[75], chanx_right_in[18], chanx_right_in[61], chany_bottom_in[1], chany_bottom_in[18], chany_bottom_in[61], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_14_sram_inv[0:3]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_7 (
		.in({chany_top_in[20], chany_top_in[62], chany_top_in[71], chanx_right_in[20], chanx_right_in[62], chany_bottom_in[2], chany_bottom_in[20], chany_bottom_in[62], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_15_sram_inv[0:3]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_9 (
		.in({chany_top_in[21], chany_top_in[64], chany_top_in[67], chanx_right_in[21], chanx_right_in[64], chany_bottom_in[3], chany_bottom_in[21], chany_bottom_in[64], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_16_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_11 (
		.in({chany_top_in[22], chany_top_in[63], chany_top_in[65], chanx_right_in[22], chanx_right_in[65], chany_bottom_in[4], chany_bottom_in[22], chany_bottom_in[65], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_17_sram_inv[0:3]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_13 (
		.in({chany_top_in[24], chany_top_in[59], chany_top_in[66], chanx_right_in[24], chanx_right_in[66], chany_bottom_in[5], chany_bottom_in[24], chany_bottom_in[66], left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_18_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_15 (
		.in({chany_top_in[25], chany_top_in[55], chany_top_in[68], chanx_right_in[25], chanx_right_in[68], chany_bottom_in[6], chany_bottom_in[25], chany_bottom_in[68], left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_19_sram_inv[0:3]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_17 (
		.in({chany_top_in[26], chany_top_in[51], chany_top_in[69], chanx_right_in[26], chanx_right_in[69], chany_bottom_in[7], chany_bottom_in[26], chany_bottom_in[69], left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_20_sram_inv[0:3]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_19 (
		.in({chany_top_in[28], chany_top_in[47], chany_top_in[70], chanx_right_in[28], chanx_right_in[70], chany_bottom_in[8], chany_bottom_in[28], chany_bottom_in[70], left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_21_sram_inv[0:3]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_21 (
		.in({chany_top_in[29], chany_top_in[43], chany_top_in[72], chanx_right_in[29], chanx_right_in[72], chany_bottom_in[9], chany_bottom_in[29], chany_bottom_in[72], left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_22_sram_inv[0:3]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_L1SB_size12 mux_left_track_23 (
		.in({chany_top_in[30], chany_top_in[39], chany_top_in[73], chanx_right_in[30], chanx_right_in[73], chany_bottom_in[10], chany_bottom_in[30], chany_bottom_in[73], left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size12_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size12_23_sram_inv[0:3]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_0 (
		.bl({bl[20:21], bl[0:1]}),
		.wl({wl[4], wl[4:5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_2 (
		.bl(bl[2:5]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_4 (
		.bl(bl[6:9]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_6 (
		.bl(bl[10:13]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_8 (
		.bl(bl[14:17]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_10 (
		.bl(bl[18:21]),
		.wl({wl[5], wl[5], wl[5], wl[5]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_12 (
		.bl(bl[0:3]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_14 (
		.bl(bl[4:7]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_16 (
		.bl(bl[8:11]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_18 (
		.bl(bl[12:15]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_20 (
		.bl(bl[16:19]),
		.wl({wl[6], wl[6], wl[6], wl[6]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_right_track_22 (
		.bl({bl[20:21], bl[0:1]}),
		.wl({wl[6], wl[6:7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_1 (
		.bl(bl[14:17]),
		.wl({wl[15], wl[15], wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_3 (
		.bl(bl[18:21]),
		.wl({wl[15], wl[15], wl[15], wl[15]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_5 (
		.bl(bl[0:3]),
		.wl({wl[16], wl[16], wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_7 (
		.bl(bl[4:7]),
		.wl({wl[16], wl[16], wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_15_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_9 (
		.bl(bl[8:11]),
		.wl({wl[16], wl[16], wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_16_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_11 (
		.bl(bl[12:15]),
		.wl({wl[16], wl[16], wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_17_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_13 (
		.bl(bl[16:19]),
		.wl({wl[16], wl[16], wl[16], wl[16]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_18_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_15 (
		.bl({bl[20:21], bl[0:1]}),
		.wl({wl[16], wl[16:17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_19_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_17 (
		.bl(bl[2:5]),
		.wl({wl[17], wl[17], wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_20_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_19 (
		.bl(bl[6:9]),
		.wl({wl[17], wl[17], wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_21_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_21 (
		.bl(bl[10:13]),
		.wl({wl[17], wl[17], wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_22_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size12_mem mem_left_track_23 (
		.bl(bl[14:17]),
		.wl({wl[17], wl[17], wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L1SB_size12_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size12_23_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size11 mux_right_track_24 (
		.in({chany_top_in[11], chany_top_in[32], chany_top_in[74], right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, chany_bottom_in[27], chany_bottom_in[32], chany_bottom_in[74], chanx_left_in[32], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L1SB_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size11_0_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_L1SB_size11 mux_right_track_26 (
		.in({chany_top_in[12], chany_top_in[33], chany_top_in[76], right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, chany_bottom_in[23], chany_bottom_in[33], chany_bottom_in[76], chanx_left_in[33], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size11_1_sram_inv[0:3]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_L1SB_size11 mux_right_track_28 (
		.in({chany_top_in[13], chany_top_in[34], chany_top_in[77], right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, chany_bottom_in[19], chany_bottom_in[34], chany_bottom_in[77], chanx_left_in[34], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size11_2_sram_inv[0:3]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_L1SB_size11 mux_right_track_30 (
		.in({chany_top_in[14], chany_top_in[36], chany_top_in[78], right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, chany_bottom_in[15], chany_bottom_in[36], chany_bottom_in[78], chanx_left_in[36], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L1SB_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size11_3_sram_inv[0:3]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_L1SB_size11 mux_left_track_25 (
		.in({chany_top_in[32], chany_top_in[35], chany_top_in[74], chanx_right_in[32], chanx_right_in[74], chany_bottom_in[11], chany_bottom_in[32], chany_bottom_in[74], left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size11_4_sram_inv[0:3]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_L1SB_size11 mux_left_track_27 (
		.in({chany_top_in[31], chany_top_in[33], chany_top_in[76], chanx_right_in[33], chanx_right_in[76], chany_bottom_in[12], chany_bottom_in[33], chany_bottom_in[76], left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size11_5_sram_inv[0:3]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_L1SB_size11 mux_left_track_29 (
		.in({chany_top_in[27], chany_top_in[34], chany_top_in[77], chanx_right_in[34], chanx_right_in[77], chany_bottom_in[13], chany_bottom_in[34], chany_bottom_in[77], left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size11_6_sram_inv[0:3]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_L1SB_size11 mux_left_track_31 (
		.in({chany_top_in[23], chany_top_in[36], chany_top_in[78], chanx_right_in[36], chanx_right_in[78], chany_bottom_in[14], chany_bottom_in[36], chany_bottom_in[78], left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size11_7_sram_inv[0:3]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_L1SB_size11_mem mem_right_track_24 (
		.bl(bl[2:5]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size11_mem mem_right_track_26 (
		.bl(bl[6:9]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size11_mem mem_right_track_28 (
		.bl(bl[10:13]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size11_mem mem_right_track_30 (
		.bl(bl[14:17]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L1SB_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size11_mem mem_left_track_25 (
		.bl(bl[18:21]),
		.wl({wl[17], wl[17], wl[17], wl[17]}),
		.mem_out(mux_tree_tapbuf_L1SB_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size11_mem mem_left_track_27 (
		.bl(bl[0:3]),
		.wl({wl[18], wl[18], wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L1SB_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size11_mem mem_left_track_29 (
		.bl(bl[4:7]),
		.wl({wl[18], wl[18], wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L1SB_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size11_mem mem_left_track_31 (
		.bl(bl[8:11]),
		.wl({wl[18], wl[18], wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L1SB_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13 mux_right_track_32 (
		.in({chany_top_in[15], chany_top_in[37], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, chany_bottom_in[14], chany_bottom_in[37], chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_0_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_L4SB_size13 mux_right_track_40 (
		.in({chany_top_in[19], chany_top_in[38], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, chany_bottom_in[13], chany_bottom_in[38], chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_1_sram_inv[0:3]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_L4SB_size13 mux_right_track_48 (
		.in({chany_top_in[23], chany_top_in[40], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_, chany_bottom_in[12], chany_bottom_in[40], chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_2_sram_inv[0:3]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_L4SB_size13 mux_right_track_56 (
		.in({chany_top_in[27], chany_top_in[41], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_, chany_bottom_in[11], chany_bottom_in[41], chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_3_sram_inv[0:3]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_L4SB_size13 mux_right_track_96 (
		.in({chany_top_in[47:48], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, chany_bottom_in[6], chany_bottom_in[48], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_4_sram_inv[0:3]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_L4SB_size13 mux_right_track_104 (
		.in({chany_top_in[49], chany_top_in[51], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, chany_bottom_in[5], chany_bottom_in[49], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size13_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_5_sram_inv[0:3]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_L4SB_size13 mux_right_track_112 (
		.in({chany_top_in[50], chany_top_in[55], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_, chany_bottom_in[4], chany_bottom_in[50], chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size13_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_6_sram_inv[0:3]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_L4SB_size13 mux_right_track_120 (
		.in({chany_top_in[52], chany_top_in[59], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_, chany_bottom_in[3], chany_bottom_in[52], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size13_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_7_sram_inv[0:3]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_33 (
		.in({chany_top_in[19], chany_top_in[37], chanx_right_in[37], chany_bottom_in[15], chany_bottom_in[37], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_8_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_41 (
		.in({chany_top_in[15], chany_top_in[38], chanx_right_in[38], chany_bottom_in[19], chany_bottom_in[38], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_9_sram_inv[0:3]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_49 (
		.in({chany_top_in[14], chany_top_in[40], chanx_right_in[40], chany_bottom_in[23], chany_bottom_in[40], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_10_sram_inv[0:3]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_57 (
		.in({chany_top_in[13], chany_top_in[41], chanx_right_in[41], chany_bottom_in[27], chany_bottom_in[41], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_11_sram_inv[0:3]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_97 (
		.in({chany_top_in[8], chany_top_in[48], chanx_right_in[48], chany_bottom_in[47:48], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_12_sram_inv[0:3]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_105 (
		.in({chany_top_in[7], chany_top_in[49], chanx_right_in[49], chany_bottom_in[49], chany_bottom_in[51], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_13_sram_inv[0:3]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_113 (
		.in({chany_top_in[6], chany_top_in[50], chanx_right_in[50], chany_bottom_in[50], chany_bottom_in[55], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_14_sram_inv[0:3]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_121 (
		.in({chany_top_in[5], chany_top_in[52], chanx_right_in[52], chany_bottom_in[52], chany_bottom_in[59], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_15_sram_inv[0:3]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_L4SB_size13_mem mem_right_track_32 (
		.bl(bl[18:21]),
		.wl({wl[7], wl[7], wl[7], wl[7]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_right_track_40 (
		.bl(bl[0:3]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_right_track_48 (
		.bl(bl[4:7]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_right_track_56 (
		.bl(bl[8:11]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_right_track_96 (
		.bl(bl[6:9]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_right_track_104 (
		.bl(bl[10:13]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_right_track_112 (
		.bl(bl[14:17]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_right_track_120 (
		.bl(bl[18:21]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_33 (
		.bl(bl[12:15]),
		.wl({wl[18], wl[18], wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_41 (
		.bl(bl[16:19]),
		.wl({wl[18], wl[18], wl[18], wl[18]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_49 (
		.bl({bl[20:21], bl[0:1]}),
		.wl({wl[18], wl[18:19], wl[19]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_57 (
		.bl(bl[2:5]),
		.wl({wl[19], wl[19], wl[19], wl[19]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_97 (
		.bl(bl[0:3]),
		.wl({wl[20], wl[20], wl[20], wl[20]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_105 (
		.bl(bl[4:7]),
		.wl({wl[20], wl[20], wl[20], wl[20]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_113 (
		.bl(bl[8:11]),
		.wl({wl[20], wl[20], wl[20], wl[20]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_121 (
		.bl(bl[12:15]),
		.wl({wl[20], wl[20], wl[20], wl[20]}),
		.mem_out(mux_tree_tapbuf_L4SB_size13_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_15_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12 mux_right_track_64 (
		.in({chany_top_in[31], chany_top_in[42], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, chany_bottom_in[10], chany_bottom_in[42], chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_0_sram_inv[0:3]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_L4SB_size12 mux_right_track_72 (
		.in({chany_top_in[35], chany_top_in[44], right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, chany_bottom_in[9], chany_bottom_in[44], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_1_sram_inv[0:3]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_L4SB_size12 mux_right_track_80 (
		.in({chany_top_in[39], chany_top_in[45], right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, chany_bottom_in[8], chany_bottom_in[45], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_2_sram_inv[0:3]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_L4SB_size12 mux_right_track_88 (
		.in({chany_top_in[43], chany_top_in[46], right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, chany_bottom_in[7], chany_bottom_in[46], chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_3_sram_inv[0:3]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_L4SB_size12 mux_right_track_128 (
		.in({chany_top_in[53], chany_top_in[63], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, chany_bottom_in[2], chany_bottom_in[53], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_4_sram_inv[0:3]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_L4SB_size12 mux_right_track_136 (
		.in({chany_top_in[54], chany_top_in[67], right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, chany_bottom_in[1], chany_bottom_in[54], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_5_sram_inv[0:3]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_L4SB_size12 mux_right_track_144 (
		.in({chany_top_in[56], chany_top_in[71], right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, chany_bottom_in[0], chany_bottom_in[56], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_6_sram_inv[0:3]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_L4SB_size12 mux_right_track_152 (
		.in({chany_top_in[57], chany_top_in[75], right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, chany_bottom_in[57], chany_bottom_in[79], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_7_sram_inv[0:3]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_65 (
		.in({chany_top_in[12], chany_top_in[42], chanx_right_in[42], chany_bottom_in[31], chany_bottom_in[42], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_8_sram_inv[0:3]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_73 (
		.in({chany_top_in[11], chany_top_in[44], chanx_right_in[44], chany_bottom_in[35], chany_bottom_in[44], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_9_sram_inv[0:3]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_81 (
		.in({chany_top_in[10], chany_top_in[45], chanx_right_in[45], chany_bottom_in[39], chany_bottom_in[45], left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_10_sram_inv[0:3]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_89 (
		.in({chany_top_in[9], chany_top_in[46], chanx_right_in[46], chany_bottom_in[43], chany_bottom_in[46], left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_11_sram_inv[0:3]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_129 (
		.in({chany_top_in[4], chany_top_in[53], chanx_right_in[53], chany_bottom_in[53], chany_bottom_in[63], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_12_sram_inv[0:3]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_137 (
		.in({chany_top_in[3], chany_top_in[54], chanx_right_in[54], chany_bottom_in[54], chany_bottom_in[67], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_13_sram_inv[0:3]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_145 (
		.in({chany_top_in[2], chany_top_in[56], chanx_right_in[56], chany_bottom_in[56], chany_bottom_in[71], left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_14_sram_inv[0:3]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_153 (
		.in({chany_top_in[1], chany_top_in[57], chanx_right_in[57], chany_bottom_in[57], chany_bottom_in[75], left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_15_sram_inv[0:3]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_L4SB_size12_mem mem_right_track_64 (
		.bl(bl[12:15]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_right_track_72 (
		.bl(bl[16:19]),
		.wl({wl[8], wl[8], wl[8], wl[8]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_right_track_80 (
		.bl({bl[20:21], bl[0:1]}),
		.wl({wl[8], wl[8:9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_right_track_88 (
		.bl(bl[2:5]),
		.wl({wl[9], wl[9], wl[9], wl[9]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_right_track_128 (
		.bl(bl[0:3]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_right_track_136 (
		.bl(bl[4:7]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_right_track_144 (
		.bl(bl[8:11]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_right_track_152 (
		.bl(bl[12:15]),
		.wl({wl[10], wl[10], wl[10], wl[10]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_65 (
		.bl(bl[6:9]),
		.wl({wl[19], wl[19], wl[19], wl[19]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_73 (
		.bl(bl[10:13]),
		.wl({wl[19], wl[19], wl[19], wl[19]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_81 (
		.bl(bl[14:17]),
		.wl({wl[19], wl[19], wl[19], wl[19]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_89 (
		.bl(bl[18:21]),
		.wl({wl[19], wl[19], wl[19], wl[19]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_129 (
		.bl(bl[16:19]),
		.wl({wl[20], wl[20], wl[20], wl[20]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_137 (
		.bl({bl[20:21], bl[0:1]}),
		.wl({wl[20], wl[20:21], wl[21]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_145 (
		.bl(bl[2:5]),
		.wl({wl[21], wl[21], wl[21], wl[21]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_153 (
		.bl(bl[6:9]),
		.wl({wl[21], wl[21], wl[21], wl[21]}),
		.mem_out(mux_tree_tapbuf_L4SB_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_15_sram_inv[0:3]));

endmodule
// ----- END Verilog module for sb_1__1_ -----

//----- Default net type -----
`default_nettype none



